module IDecode(
  input         clock,
  input         reset,
  input         io_rst_n,
  input  [31:0] io_pc_i,
  input  [31:0] io_inst_i,
  input  [31:0] io_excepttype_i,
  input         io_not_stall_i,
  input  [7:0]  io_ex_aluop_i,
  input         io_ex_wreg_i,
  input  [31:0] io_ex_wdata_i,
  input  [4:0]  io_ex_wd_i,
  input         io_mem_wreg_i,
  input  [31:0] io_mem_wdata_i,
  input  [4:0]  io_mem_wd_i,
  input         io_ex_csr_reg_we_i,
  input         io_mem_csr_reg_we_i,
  input         io_wb_csr_reg_we_i,
  input         io_ex_not_stall_i,
  input         io_mem_not_stall_i,
  input  [31:0] io_reg1_data_i,
  input  [31:0] io_reg2_data_i,
  input         io_is_in_delayslot_i,
  input         io_step_i,
  input  [1:0]  io_prv_i,
  input  [31:0] io_csr_reg_data_i,
  input         io_csr_protect_i,
  output [31:0] io_csr_reg_data_o,
  output        io_csr_reg_read_o,
  output        io_csr_reg_we_o,
  output [11:0] io_csr_reg_addr_o,
  output        io_reg1_read_o,
  output        io_reg2_read_o,
  output [4:0]  io_reg1_addr_o,
  output [4:0]  io_reg2_addr_o,
  output [7:0]  io_aluop_o,
  output [2:0]  io_alusel_o,
  output [31:0] io_reg1_o,
  output [31:0] io_reg2_o,
  output [31:0] io_mem_addr_o,
  output [4:0]  io_wd_o,
  output        io_wreg_o,
  output [31:0] io_inst_o,
  output        io_next_inst_in_delayslot_o,
  output        io_branch_flag_o,
  output [31:0] io_branch_target_address_o,
  output [31:0] io_link_addr_o,
  output        io_is_in_delayslot_o,
  output [31:0] io_excepttype_o,
  output [31:0] io_current_inst_address_o,
  output        io_not_stall_o,
  output        io_step_o,
  output        io_stallreq
);
  reg [31:0] imm; // @[IDecode.scala 203:15]
  reg [31:0] _RAND_0;
  reg [31:0] imm_i_type; // @[IDecode.scala 204:22]
  reg [31:0] _RAND_1;
  reg [31:0] imm_s_type; // @[IDecode.scala 205:22]
  reg [31:0] _RAND_2;
  reg [31:0] imm_u_type; // @[IDecode.scala 206:22]
  reg [31:0] _RAND_3;
  reg [31:0] imm_sb_type; // @[IDecode.scala 207:23]
  reg [31:0] _RAND_4;
  reg [31:0] imm_uj_type; // @[IDecode.scala 208:23]
  reg [31:0] _RAND_5;
  reg [31:0] zimm; // @[IDecode.scala 209:16]
  reg [31:0] _RAND_6;
  wire [19:0] _T_12; // @[Bitwise.scala 71:12]
  wire [26:0] _T_19; // @[Cat.scala 29:58]
  wire [18:0] _T_27; // @[Bitwise.scala 71:12]
  wire [30:0] _T_35; // @[Cat.scala 29:58]
  wire [10:0] _T_39; // @[Bitwise.scala 71:12]
  wire [30:0] _T_47; // @[Cat.scala 29:58]
  reg  instvalid; // @[IDecode.scala 219:21]
  reg [31:0] _RAND_7;
  reg  stallreq_for_reg1_loadrelate; // @[IDecode.scala 221:40]
  reg [31:0] _RAND_8;
  reg  stallreq_for_reg2_loadrelate; // @[IDecode.scala 222:40]
  reg [31:0] _RAND_9;
  reg  stallreq_for_csr_write_relate; // @[IDecode.scala 224:41]
  reg [31:0] _RAND_10;
  reg  stallreq_for_csr_read_relate; // @[IDecode.scala 225:40]
  reg [31:0] _RAND_11;
  reg  pre_inst_is_load; // @[IDecode.scala 226:28]
  reg [31:0] _RAND_12;
  reg  excepttype_is_syscall; // @[IDecode.scala 227:33]
  reg [31:0] _RAND_13;
  reg  excepttype_is_break; // @[IDecode.scala 228:31]
  reg [31:0] _RAND_14;
  reg  excepttype_is_sret; // @[IDecode.scala 229:30]
  reg [31:0] _RAND_15;
  reg  excepttype_is_mret; // @[IDecode.scala 230:30]
  reg [31:0] _RAND_16;
  reg  excepttype_is_fence_i; // @[IDecode.scala 231:33]
  reg [31:0] _RAND_17;
  wire  _T_54; // @[IDecode.scala 236:44]
  wire  _T_56; // @[IDecode.scala 236:89]
  wire  _T_59; // @[IDecode.scala 239:94]
  wire  _T_61; // @[IDecode.scala 241:46]
  wire  _T_62; // @[IDecode.scala 241:77]
  wire  _T_64; // @[IDecode.scala 244:20]
  wire  _T_65; // @[IDecode.scala 244:55]
  wire  _T_66; // @[IDecode.scala 244:37]
  wire  _T_67; // @[IDecode.scala 244:91]
  wire  _T_68; // @[IDecode.scala 244:73]
  wire  _T_69; // @[IDecode.scala 245:20]
  wire  _T_70; // @[IDecode.scala 244:108]
  wire  _T_71; // @[IDecode.scala 245:56]
  wire  _T_72; // @[IDecode.scala 245:38]
  wire  _T_73; // @[IDecode.scala 245:91]
  wire  _T_74; // @[IDecode.scala 245:73]
  wire  _T_75; // @[IDecode.scala 246:20]
  wire  _T_76; // @[IDecode.scala 245:108]
  wire  _T_77; // @[IDecode.scala 246:55]
  wire  _T_78; // @[IDecode.scala 246:37]
  wire  _T_79; // @[IDecode.scala 246:97]
  wire  _T_80; // @[IDecode.scala 246:79]
  wire  _T_81; // @[IDecode.scala 247:20]
  wire  _T_82; // @[IDecode.scala 246:120]
  wire  _T_83; // @[IDecode.scala 247:61]
  wire  _T_84; // @[IDecode.scala 247:43]
  wire  _T_85; // @[IDecode.scala 247:102]
  wire  _T_86; // @[IDecode.scala 247:84]
  wire  _T_87; // @[IDecode.scala 248:20]
  wire  _T_88; // @[IDecode.scala 247:124]
  wire  _T_89; // @[IDecode.scala 248:61]
  wire  _T_90; // @[IDecode.scala 248:43]
  wire  _T_91; // @[IDecode.scala 248:102]
  wire  _T_92; // @[IDecode.scala 248:84]
  wire  _T_93; // @[IDecode.scala 249:20]
  wire  _T_130; // @[IDecode.scala 265:56]
  wire  _T_131; // @[Conditional.scala 37:30]
  wire  _T_132; // @[Conditional.scala 37:30]
  wire  _T_133; // @[Conditional.scala 37:30]
  wire  _GEN_0; // @[Conditional.scala 39:67]
  wire  _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_2; // @[Conditional.scala 39:67]
  wire  _GEN_3; // @[Conditional.scala 40:58]
  wire  _GEN_4; // @[Conditional.scala 40:58]
  wire  _GEN_5; // @[Conditional.scala 40:58]
  wire  _GEN_8; // @[IDecode.scala 259:52]
  wire  excepttype_b_1; // @[IDecode.scala 256:32]
  wire  _GEN_7; // @[IDecode.scala 259:52]
  wire  excepttype_b_0; // @[IDecode.scala 256:32]
  wire  _GEN_10; // @[IDecode.scala 259:52]
  wire  excepttype_b_3; // @[IDecode.scala 256:32]
  wire  _GEN_9; // @[IDecode.scala 259:52]
  wire  excepttype_b_2; // @[IDecode.scala 256:32]
  wire  _GEN_12; // @[IDecode.scala 259:52]
  wire  excepttype_b_5; // @[IDecode.scala 256:32]
  wire  _GEN_11; // @[IDecode.scala 259:52]
  wire  excepttype_b_4; // @[IDecode.scala 256:32]
  wire  _GEN_14; // @[IDecode.scala 259:52]
  wire  excepttype_b_7; // @[IDecode.scala 256:32]
  wire  _GEN_13; // @[IDecode.scala 259:52]
  wire  excepttype_b_6; // @[IDecode.scala 256:32]
  wire [7:0] _T_140; // @[IDecode.scala 278:35]
  wire  _GEN_16; // @[IDecode.scala 259:52]
  wire  excepttype_b_9; // @[IDecode.scala 256:32]
  wire  _GEN_15; // @[IDecode.scala 259:52]
  wire  excepttype_b_8; // @[IDecode.scala 256:32]
  wire  _GEN_18; // @[IDecode.scala 259:52]
  wire  excepttype_b_11; // @[IDecode.scala 256:32]
  wire  _GEN_17; // @[IDecode.scala 259:52]
  wire  excepttype_b_10; // @[IDecode.scala 256:32]
  wire  _GEN_20; // @[IDecode.scala 259:52]
  wire  excepttype_b_13; // @[IDecode.scala 256:32]
  wire  _GEN_19; // @[IDecode.scala 259:52]
  wire  excepttype_b_12; // @[IDecode.scala 256:32]
  wire  _GEN_22; // @[IDecode.scala 259:52]
  wire  excepttype_b_15; // @[IDecode.scala 256:32]
  wire  _GEN_21; // @[IDecode.scala 259:52]
  wire  excepttype_b_14; // @[IDecode.scala 256:32]
  wire [15:0] _T_148; // @[IDecode.scala 278:35]
  wire  _GEN_24; // @[IDecode.scala 259:52]
  wire  excepttype_b_17; // @[IDecode.scala 256:32]
  wire  _GEN_23; // @[IDecode.scala 259:52]
  wire  excepttype_b_16; // @[IDecode.scala 256:32]
  wire  _GEN_26; // @[IDecode.scala 259:52]
  wire  excepttype_b_19; // @[IDecode.scala 256:32]
  wire  _GEN_25; // @[IDecode.scala 259:52]
  wire  excepttype_b_18; // @[IDecode.scala 256:32]
  wire  _GEN_28; // @[IDecode.scala 259:52]
  wire  excepttype_b_21; // @[IDecode.scala 256:32]
  wire  _GEN_27; // @[IDecode.scala 259:52]
  wire  excepttype_b_20; // @[IDecode.scala 256:32]
  wire  _GEN_30; // @[IDecode.scala 259:52]
  wire  excepttype_b_23; // @[IDecode.scala 256:32]
  wire  _GEN_29; // @[IDecode.scala 259:52]
  wire  excepttype_b_22; // @[IDecode.scala 256:32]
  wire [7:0] _T_155; // @[IDecode.scala 278:35]
  wire  _GEN_32; // @[IDecode.scala 259:52]
  wire  excepttype_b_25; // @[IDecode.scala 256:32]
  wire  _GEN_31; // @[IDecode.scala 259:52]
  wire  excepttype_b_24; // @[IDecode.scala 256:32]
  wire  _GEN_34; // @[IDecode.scala 259:52]
  wire  excepttype_b_27; // @[IDecode.scala 256:32]
  wire  _GEN_33; // @[IDecode.scala 259:52]
  wire  excepttype_b_26; // @[IDecode.scala 256:32]
  wire  _GEN_36; // @[IDecode.scala 259:52]
  wire  excepttype_b_29; // @[IDecode.scala 256:32]
  wire  _GEN_35; // @[IDecode.scala 259:52]
  wire  excepttype_b_28; // @[IDecode.scala 256:32]
  wire  _GEN_38; // @[IDecode.scala 259:52]
  wire  excepttype_b_31; // @[IDecode.scala 256:32]
  wire  _GEN_37; // @[IDecode.scala 259:52]
  wire  excepttype_b_30; // @[IDecode.scala 256:32]
  wire [31:0] _T_164; // @[IDecode.scala 278:35]
  wire  _GEN_6; // @[IDecode.scala 259:52]
  wire [31:0] _GEN_39; // @[IDecode.scala 259:52]
  wire  _T_167; // @[IDecode.scala 285:32]
  wire  _T_168; // @[IDecode.scala 285:93]
  wire  _T_170; // @[IDecode.scala 285:74]
  wire [31:0] _T_172; // @[IDecode.scala 444:19]
  wire [31:0] _T_174; // @[IDecode.scala 620:16]
  wire [31:0] _T_176; // @[IDecode.scala 629:32]
  wire [31:0] _T_178; // @[Cat.scala 29:58]
  wire  _T_179; // @[IDecode.scala 639:23]
  wire [31:0] _T_181; // @[IDecode.scala 639:46]
  wire [31:0] _T_182; // @[IDecode.scala 639:12]
  wire  _T_187; // @[IDecode.scala 648:23]
  wire [31:0] _T_190; // @[IDecode.scala 648:12]
  wire  _T_197; // @[IDecode.scala 657:30]
  wire [31:0] _T_200; // @[IDecode.scala 657:12]
  wire  _T_209; // @[IDecode.scala 666:23]
  wire [31:0] _T_212; // @[IDecode.scala 666:12]
  wire  _T_219; // @[IDecode.scala 675:30]
  wire [31:0] _T_222; // @[IDecode.scala 675:12]
  wire  _T_231; // @[IDecode.scala 684:23]
  wire [31:0] _T_234; // @[IDecode.scala 684:12]
  wire [31:0] _T_240; // @[IDecode.scala 693:21]
  wire [31:0] _T_250; // @[IDecode.scala 739:21]
  wire  _T_255; // @[IDecode.scala 764:60]
  wire  _T_256; // @[IDecode.scala 764:89]
  wire  _T_257; // @[IDecode.scala 764:78]
  wire  _T_259; // @[IDecode.scala 764:127]
  wire  _T_260; // @[IDecode.scala 764:107]
  wire  _T_265; // @[IDecode.scala 773:121]
  wire  _T_266; // @[IDecode.scala 773:107]
  wire  _T_274; // @[IDecode.scala 810:54]
  wire  _T_278; // @[IDecode.scala 835:21]
  wire  _T_280; // @[IDecode.scala 844:42]
  wire [31:0] _T_290; // @[Lookup.scala 31:38]
  wire  _T_291; // @[Lookup.scala 31:38]
  wire  _T_293; // @[Lookup.scala 31:38]
  wire  _T_295; // @[Lookup.scala 31:38]
  wire  _T_297; // @[Lookup.scala 31:38]
  wire  _T_299; // @[Lookup.scala 31:38]
  wire  _T_301; // @[Lookup.scala 31:38]
  wire [31:0] _T_302; // @[Lookup.scala 31:38]
  wire  _T_303; // @[Lookup.scala 31:38]
  wire  _T_305; // @[Lookup.scala 31:38]
  wire  _T_307; // @[Lookup.scala 31:38]
  wire [31:0] _T_308; // @[Lookup.scala 31:38]
  wire  _T_309; // @[Lookup.scala 31:38]
  wire  _T_311; // @[Lookup.scala 31:38]
  wire [31:0] _T_312; // @[Lookup.scala 31:38]
  wire  _T_313; // @[Lookup.scala 31:38]
  wire  _T_315; // @[Lookup.scala 31:38]
  wire  _T_317; // @[Lookup.scala 31:38]
  wire  _T_319; // @[Lookup.scala 31:38]
  wire  _T_321; // @[Lookup.scala 31:38]
  wire  _T_323; // @[Lookup.scala 31:38]
  wire  _T_325; // @[Lookup.scala 31:38]
  wire  _T_327; // @[Lookup.scala 31:38]
  wire  _T_329; // @[Lookup.scala 31:38]
  wire  _T_331; // @[Lookup.scala 31:38]
  wire  _T_333; // @[Lookup.scala 31:38]
  wire  _T_335; // @[Lookup.scala 31:38]
  wire  _T_337; // @[Lookup.scala 31:38]
  wire  _T_339; // @[Lookup.scala 31:38]
  wire  _T_341; // @[Lookup.scala 31:38]
  wire  _T_343; // @[Lookup.scala 31:38]
  wire  _T_345; // @[Lookup.scala 31:38]
  wire  _T_347; // @[Lookup.scala 31:38]
  wire  _T_349; // @[Lookup.scala 31:38]
  wire  _T_351; // @[Lookup.scala 31:38]
  wire  _T_353; // @[Lookup.scala 31:38]
  wire  _T_355; // @[Lookup.scala 31:38]
  wire  _T_357; // @[Lookup.scala 31:38]
  wire  _T_359; // @[Lookup.scala 31:38]
  wire  _T_361; // @[Lookup.scala 31:38]
  wire  _T_363; // @[Lookup.scala 31:38]
  wire  _T_365; // @[Lookup.scala 31:38]
  wire  _T_367; // @[Lookup.scala 31:38]
  wire  _T_369; // @[Lookup.scala 31:38]
  wire  _T_371; // @[Lookup.scala 31:38]
  wire  _T_373; // @[Lookup.scala 31:38]
  wire  _T_375; // @[Lookup.scala 31:38]
  wire  _T_377; // @[Lookup.scala 31:38]
  wire  _T_379; // @[Lookup.scala 31:38]
  wire  _T_381; // @[Lookup.scala 31:38]
  wire  _T_383; // @[Lookup.scala 31:38]
  wire  _T_385; // @[Lookup.scala 31:38]
  wire  _T_387; // @[Lookup.scala 31:38]
  wire  _T_389; // @[Lookup.scala 31:38]
  wire  _T_391; // @[Lookup.scala 31:38]
  wire  _T_393; // @[Lookup.scala 31:38]
  wire  _T_395; // @[Lookup.scala 31:38]
  wire  _T_397; // @[Lookup.scala 31:38]
  wire  _T_399; // @[Lookup.scala 31:38]
  wire  _T_401; // @[Lookup.scala 31:38]
  wire  _T_403; // @[Lookup.scala 31:38]
  wire  _T_405; // @[Lookup.scala 31:38]
  wire [31:0] _T_406; // @[Lookup.scala 31:38]
  wire  _T_407; // @[Lookup.scala 31:38]
  wire [31:0] _T_408; // @[Lookup.scala 31:38]
  wire  _T_409; // @[Lookup.scala 31:38]
  wire  _T_411; // @[Lookup.scala 31:38]
  wire  _T_413; // @[Lookup.scala 31:38]
  wire  _T_415; // @[Lookup.scala 31:38]
  wire  _T_417; // @[Lookup.scala 31:38]
  wire  _T_419; // @[Lookup.scala 31:38]
  wire  _T_421; // @[Lookup.scala 31:38]
  wire  _T_423; // @[Lookup.scala 31:38]
  wire  _T_425; // @[Lookup.scala 31:38]
  wire  _T_427; // @[Lookup.scala 31:38]
  wire [7:0] _T_428; // @[Lookup.scala 33:37]
  wire [7:0] _T_429; // @[Lookup.scala 33:37]
  wire [7:0] _T_430; // @[Lookup.scala 33:37]
  wire [7:0] _T_431; // @[Lookup.scala 33:37]
  wire [7:0] _T_432; // @[Lookup.scala 33:37]
  wire [7:0] _T_433; // @[Lookup.scala 33:37]
  wire [7:0] _T_434; // @[Lookup.scala 33:37]
  wire [7:0] _T_435; // @[Lookup.scala 33:37]
  wire [7:0] _T_436; // @[Lookup.scala 33:37]
  wire [7:0] _T_437; // @[Lookup.scala 33:37]
  wire [7:0] _T_438; // @[Lookup.scala 33:37]
  wire [7:0] _T_439; // @[Lookup.scala 33:37]
  wire [7:0] _T_440; // @[Lookup.scala 33:37]
  wire [7:0] _T_441; // @[Lookup.scala 33:37]
  wire [7:0] _T_442; // @[Lookup.scala 33:37]
  wire [7:0] _T_443; // @[Lookup.scala 33:37]
  wire [7:0] _T_444; // @[Lookup.scala 33:37]
  wire [7:0] _T_445; // @[Lookup.scala 33:37]
  wire [7:0] _T_446; // @[Lookup.scala 33:37]
  wire [7:0] _T_447; // @[Lookup.scala 33:37]
  wire [7:0] _T_448; // @[Lookup.scala 33:37]
  wire [7:0] _T_449; // @[Lookup.scala 33:37]
  wire [7:0] _T_450; // @[Lookup.scala 33:37]
  wire [7:0] _T_451; // @[Lookup.scala 33:37]
  wire [7:0] _T_452; // @[Lookup.scala 33:37]
  wire [7:0] _T_453; // @[Lookup.scala 33:37]
  wire [7:0] _T_454; // @[Lookup.scala 33:37]
  wire [7:0] _T_455; // @[Lookup.scala 33:37]
  wire [7:0] _T_456; // @[Lookup.scala 33:37]
  wire [7:0] _T_457; // @[Lookup.scala 33:37]
  wire [7:0] _T_458; // @[Lookup.scala 33:37]
  wire [7:0] _T_459; // @[Lookup.scala 33:37]
  wire [7:0] _T_460; // @[Lookup.scala 33:37]
  wire [7:0] _T_461; // @[Lookup.scala 33:37]
  wire [7:0] _T_462; // @[Lookup.scala 33:37]
  wire [7:0] _T_463; // @[Lookup.scala 33:37]
  wire [7:0] _T_464; // @[Lookup.scala 33:37]
  wire [7:0] _T_465; // @[Lookup.scala 33:37]
  wire [7:0] _T_466; // @[Lookup.scala 33:37]
  wire [7:0] _T_467; // @[Lookup.scala 33:37]
  wire [7:0] _T_468; // @[Lookup.scala 33:37]
  wire [7:0] _T_469; // @[Lookup.scala 33:37]
  wire [7:0] _T_470; // @[Lookup.scala 33:37]
  wire [7:0] _T_471; // @[Lookup.scala 33:37]
  wire [7:0] _T_472; // @[Lookup.scala 33:37]
  wire [7:0] _T_473; // @[Lookup.scala 33:37]
  wire [7:0] _T_474; // @[Lookup.scala 33:37]
  wire [7:0] _T_475; // @[Lookup.scala 33:37]
  wire [7:0] _T_476; // @[Lookup.scala 33:37]
  wire [7:0] _T_477; // @[Lookup.scala 33:37]
  wire [7:0] _T_478; // @[Lookup.scala 33:37]
  wire [7:0] _T_479; // @[Lookup.scala 33:37]
  wire [7:0] _T_480; // @[Lookup.scala 33:37]
  wire [7:0] _T_481; // @[Lookup.scala 33:37]
  wire [7:0] _T_482; // @[Lookup.scala 33:37]
  wire [7:0] _T_483; // @[Lookup.scala 33:37]
  wire [7:0] _T_484; // @[Lookup.scala 33:37]
  wire [7:0] _T_485; // @[Lookup.scala 33:37]
  wire [7:0] _T_486; // @[Lookup.scala 33:37]
  wire [7:0] _T_487; // @[Lookup.scala 33:37]
  wire [7:0] _T_488; // @[Lookup.scala 33:37]
  wire [7:0] _T_489; // @[Lookup.scala 33:37]
  wire [7:0] _T_490; // @[Lookup.scala 33:37]
  wire [7:0] _T_491; // @[Lookup.scala 33:37]
  wire [7:0] _T_492; // @[Lookup.scala 33:37]
  wire [7:0] _T_493; // @[Lookup.scala 33:37]
  wire [7:0] _T_494; // @[Lookup.scala 33:37]
  wire [7:0] _T_495; // @[Lookup.scala 33:37]
  wire [7:0] _T_496; // @[Lookup.scala 33:37]
  wire [2:0] _T_497; // @[Lookup.scala 33:37]
  wire [2:0] _T_498; // @[Lookup.scala 33:37]
  wire [2:0] _T_499; // @[Lookup.scala 33:37]
  wire [2:0] _T_500; // @[Lookup.scala 33:37]
  wire [2:0] _T_501; // @[Lookup.scala 33:37]
  wire [2:0] _T_502; // @[Lookup.scala 33:37]
  wire [2:0] _T_503; // @[Lookup.scala 33:37]
  wire [2:0] _T_504; // @[Lookup.scala 33:37]
  wire [2:0] _T_505; // @[Lookup.scala 33:37]
  wire [2:0] _T_506; // @[Lookup.scala 33:37]
  wire [2:0] _T_507; // @[Lookup.scala 33:37]
  wire [2:0] _T_508; // @[Lookup.scala 33:37]
  wire [2:0] _T_509; // @[Lookup.scala 33:37]
  wire [2:0] _T_510; // @[Lookup.scala 33:37]
  wire [2:0] _T_511; // @[Lookup.scala 33:37]
  wire [2:0] _T_512; // @[Lookup.scala 33:37]
  wire [2:0] _T_513; // @[Lookup.scala 33:37]
  wire [2:0] _T_514; // @[Lookup.scala 33:37]
  wire [2:0] _T_515; // @[Lookup.scala 33:37]
  wire [2:0] _T_516; // @[Lookup.scala 33:37]
  wire [2:0] _T_517; // @[Lookup.scala 33:37]
  wire [2:0] _T_518; // @[Lookup.scala 33:37]
  wire [2:0] _T_519; // @[Lookup.scala 33:37]
  wire [2:0] _T_520; // @[Lookup.scala 33:37]
  wire [2:0] _T_521; // @[Lookup.scala 33:37]
  wire [2:0] _T_522; // @[Lookup.scala 33:37]
  wire [2:0] _T_523; // @[Lookup.scala 33:37]
  wire [2:0] _T_524; // @[Lookup.scala 33:37]
  wire [2:0] _T_525; // @[Lookup.scala 33:37]
  wire [2:0] _T_526; // @[Lookup.scala 33:37]
  wire [2:0] _T_527; // @[Lookup.scala 33:37]
  wire [2:0] _T_528; // @[Lookup.scala 33:37]
  wire [2:0] _T_529; // @[Lookup.scala 33:37]
  wire [2:0] _T_530; // @[Lookup.scala 33:37]
  wire [2:0] _T_531; // @[Lookup.scala 33:37]
  wire [2:0] _T_532; // @[Lookup.scala 33:37]
  wire [2:0] _T_533; // @[Lookup.scala 33:37]
  wire [2:0] _T_534; // @[Lookup.scala 33:37]
  wire [2:0] _T_535; // @[Lookup.scala 33:37]
  wire [2:0] _T_536; // @[Lookup.scala 33:37]
  wire [2:0] _T_537; // @[Lookup.scala 33:37]
  wire [2:0] _T_538; // @[Lookup.scala 33:37]
  wire [2:0] _T_539; // @[Lookup.scala 33:37]
  wire [2:0] _T_540; // @[Lookup.scala 33:37]
  wire [2:0] _T_541; // @[Lookup.scala 33:37]
  wire [2:0] _T_542; // @[Lookup.scala 33:37]
  wire [2:0] _T_543; // @[Lookup.scala 33:37]
  wire [2:0] _T_544; // @[Lookup.scala 33:37]
  wire [2:0] _T_545; // @[Lookup.scala 33:37]
  wire [2:0] _T_546; // @[Lookup.scala 33:37]
  wire [2:0] _T_547; // @[Lookup.scala 33:37]
  wire [2:0] _T_548; // @[Lookup.scala 33:37]
  wire [2:0] _T_549; // @[Lookup.scala 33:37]
  wire [2:0] _T_550; // @[Lookup.scala 33:37]
  wire [2:0] _T_551; // @[Lookup.scala 33:37]
  wire [2:0] _T_552; // @[Lookup.scala 33:37]
  wire [2:0] _T_553; // @[Lookup.scala 33:37]
  wire [2:0] _T_554; // @[Lookup.scala 33:37]
  wire [2:0] _T_555; // @[Lookup.scala 33:37]
  wire [2:0] _T_556; // @[Lookup.scala 33:37]
  wire [2:0] _T_557; // @[Lookup.scala 33:37]
  wire [2:0] _T_558; // @[Lookup.scala 33:37]
  wire [2:0] _T_559; // @[Lookup.scala 33:37]
  wire [2:0] _T_560; // @[Lookup.scala 33:37]
  wire [2:0] _T_561; // @[Lookup.scala 33:37]
  wire [2:0] _T_562; // @[Lookup.scala 33:37]
  wire [2:0] _T_563; // @[Lookup.scala 33:37]
  wire [2:0] _T_564; // @[Lookup.scala 33:37]
  wire [2:0] _T_565; // @[Lookup.scala 33:37]
  wire  _T_636; // @[Lookup.scala 33:37]
  wire  _T_637; // @[Lookup.scala 33:37]
  wire  _T_638; // @[Lookup.scala 33:37]
  wire  _T_639; // @[Lookup.scala 33:37]
  wire  _T_640; // @[Lookup.scala 33:37]
  wire  _T_641; // @[Lookup.scala 33:37]
  wire  _T_642; // @[Lookup.scala 33:37]
  wire  _T_643; // @[Lookup.scala 33:37]
  wire  _T_644; // @[Lookup.scala 33:37]
  wire  _T_645; // @[Lookup.scala 33:37]
  wire  _T_646; // @[Lookup.scala 33:37]
  wire  _T_647; // @[Lookup.scala 33:37]
  wire  _T_648; // @[Lookup.scala 33:37]
  wire  _T_649; // @[Lookup.scala 33:37]
  wire  _T_650; // @[Lookup.scala 33:37]
  wire  _T_651; // @[Lookup.scala 33:37]
  wire  _T_652; // @[Lookup.scala 33:37]
  wire  _T_653; // @[Lookup.scala 33:37]
  wire  _T_654; // @[Lookup.scala 33:37]
  wire  _T_655; // @[Lookup.scala 33:37]
  wire  _T_656; // @[Lookup.scala 33:37]
  wire  _T_657; // @[Lookup.scala 33:37]
  wire  _T_658; // @[Lookup.scala 33:37]
  wire  _T_659; // @[Lookup.scala 33:37]
  wire  _T_660; // @[Lookup.scala 33:37]
  wire  _T_661; // @[Lookup.scala 33:37]
  wire  _T_662; // @[Lookup.scala 33:37]
  wire  _T_663; // @[Lookup.scala 33:37]
  wire  _T_664; // @[Lookup.scala 33:37]
  wire  _T_665; // @[Lookup.scala 33:37]
  wire  _T_666; // @[Lookup.scala 33:37]
  wire  _T_667; // @[Lookup.scala 33:37]
  wire  _T_668; // @[Lookup.scala 33:37]
  wire  _T_669; // @[Lookup.scala 33:37]
  wire  _T_670; // @[Lookup.scala 33:37]
  wire  _T_671; // @[Lookup.scala 33:37]
  wire  _T_672; // @[Lookup.scala 33:37]
  wire  _T_673; // @[Lookup.scala 33:37]
  wire  _T_674; // @[Lookup.scala 33:37]
  wire  _T_675; // @[Lookup.scala 33:37]
  wire  _T_676; // @[Lookup.scala 33:37]
  wire  _T_677; // @[Lookup.scala 33:37]
  wire  _T_678; // @[Lookup.scala 33:37]
  wire  _T_679; // @[Lookup.scala 33:37]
  wire  _T_680; // @[Lookup.scala 33:37]
  wire  _T_681; // @[Lookup.scala 33:37]
  wire  _T_682; // @[Lookup.scala 33:37]
  wire  _T_683; // @[Lookup.scala 33:37]
  wire  _T_684; // @[Lookup.scala 33:37]
  wire  _T_685; // @[Lookup.scala 33:37]
  wire  _T_686; // @[Lookup.scala 33:37]
  wire  _T_687; // @[Lookup.scala 33:37]
  wire  _T_688; // @[Lookup.scala 33:37]
  wire  _T_689; // @[Lookup.scala 33:37]
  wire  _T_690; // @[Lookup.scala 33:37]
  wire  _T_691; // @[Lookup.scala 33:37]
  wire  _T_692; // @[Lookup.scala 33:37]
  wire  _T_693; // @[Lookup.scala 33:37]
  wire  _T_694; // @[Lookup.scala 33:37]
  wire  _T_695; // @[Lookup.scala 33:37]
  wire  _T_696; // @[Lookup.scala 33:37]
  wire  _T_697; // @[Lookup.scala 33:37]
  wire  _T_698; // @[Lookup.scala 33:37]
  wire  _T_699; // @[Lookup.scala 33:37]
  wire  _T_700; // @[Lookup.scala 33:37]
  wire  _T_701; // @[Lookup.scala 33:37]
  wire  _T_702; // @[Lookup.scala 33:37]
  wire  _T_703; // @[Lookup.scala 33:37]
  wire  _T_728; // @[Lookup.scala 33:37]
  wire  _T_729; // @[Lookup.scala 33:37]
  wire  _T_730; // @[Lookup.scala 33:37]
  wire  _T_731; // @[Lookup.scala 33:37]
  wire  _T_732; // @[Lookup.scala 33:37]
  wire  _T_733; // @[Lookup.scala 33:37]
  wire  _T_734; // @[Lookup.scala 33:37]
  wire  _T_735; // @[Lookup.scala 33:37]
  wire  _T_736; // @[Lookup.scala 33:37]
  wire  _T_737; // @[Lookup.scala 33:37]
  wire  _T_738; // @[Lookup.scala 33:37]
  wire  _T_739; // @[Lookup.scala 33:37]
  wire  _T_740; // @[Lookup.scala 33:37]
  wire  _T_741; // @[Lookup.scala 33:37]
  wire  _T_742; // @[Lookup.scala 33:37]
  wire  _T_743; // @[Lookup.scala 33:37]
  wire  _T_744; // @[Lookup.scala 33:37]
  wire  _T_745; // @[Lookup.scala 33:37]
  wire  _T_746; // @[Lookup.scala 33:37]
  wire  _T_747; // @[Lookup.scala 33:37]
  wire  _T_748; // @[Lookup.scala 33:37]
  wire  _T_749; // @[Lookup.scala 33:37]
  wire  _T_750; // @[Lookup.scala 33:37]
  wire  _T_751; // @[Lookup.scala 33:37]
  wire  _T_752; // @[Lookup.scala 33:37]
  wire  _T_753; // @[Lookup.scala 33:37]
  wire  _T_754; // @[Lookup.scala 33:37]
  wire  _T_755; // @[Lookup.scala 33:37]
  wire  _T_756; // @[Lookup.scala 33:37]
  wire  _T_757; // @[Lookup.scala 33:37]
  wire  _T_758; // @[Lookup.scala 33:37]
  wire  _T_759; // @[Lookup.scala 33:37]
  wire  _T_760; // @[Lookup.scala 33:37]
  wire  _T_761; // @[Lookup.scala 33:37]
  wire  _T_762; // @[Lookup.scala 33:37]
  wire  _T_763; // @[Lookup.scala 33:37]
  wire  _T_764; // @[Lookup.scala 33:37]
  wire  _T_765; // @[Lookup.scala 33:37]
  wire  _T_766; // @[Lookup.scala 33:37]
  wire  _T_767; // @[Lookup.scala 33:37]
  wire  _T_768; // @[Lookup.scala 33:37]
  wire  _T_769; // @[Lookup.scala 33:37]
  wire  _T_770; // @[Lookup.scala 33:37]
  wire  _T_771; // @[Lookup.scala 33:37]
  wire  _T_772; // @[Lookup.scala 33:37]
  wire  _T_783; // @[Lookup.scala 33:37]
  wire  _T_784; // @[Lookup.scala 33:37]
  wire  _T_785; // @[Lookup.scala 33:37]
  wire  _T_786; // @[Lookup.scala 33:37]
  wire  _T_787; // @[Lookup.scala 33:37]
  wire  _T_788; // @[Lookup.scala 33:37]
  wire  _T_789; // @[Lookup.scala 33:37]
  wire  _T_790; // @[Lookup.scala 33:37]
  wire  _T_791; // @[Lookup.scala 33:37]
  wire  _T_792; // @[Lookup.scala 33:37]
  wire  _T_793; // @[Lookup.scala 33:37]
  wire  _T_794; // @[Lookup.scala 33:37]
  wire  _T_795; // @[Lookup.scala 33:37]
  wire  _T_796; // @[Lookup.scala 33:37]
  wire  _T_797; // @[Lookup.scala 33:37]
  wire  _T_798; // @[Lookup.scala 33:37]
  wire  _T_799; // @[Lookup.scala 33:37]
  wire  _T_800; // @[Lookup.scala 33:37]
  wire  _T_801; // @[Lookup.scala 33:37]
  wire  _T_802; // @[Lookup.scala 33:37]
  wire  _T_803; // @[Lookup.scala 33:37]
  wire  _T_804; // @[Lookup.scala 33:37]
  wire  _T_805; // @[Lookup.scala 33:37]
  wire  _T_806; // @[Lookup.scala 33:37]
  wire  _T_807; // @[Lookup.scala 33:37]
  wire  _T_808; // @[Lookup.scala 33:37]
  wire  _T_809; // @[Lookup.scala 33:37]
  wire  _T_810; // @[Lookup.scala 33:37]
  wire  _T_811; // @[Lookup.scala 33:37]
  wire  _T_812; // @[Lookup.scala 33:37]
  wire  _T_813; // @[Lookup.scala 33:37]
  wire  _T_814; // @[Lookup.scala 33:37]
  wire  _T_815; // @[Lookup.scala 33:37]
  wire  _T_816; // @[Lookup.scala 33:37]
  wire  _T_817; // @[Lookup.scala 33:37]
  wire  _T_818; // @[Lookup.scala 33:37]
  wire  _T_819; // @[Lookup.scala 33:37]
  wire  _T_820; // @[Lookup.scala 33:37]
  wire  _T_821; // @[Lookup.scala 33:37]
  wire  _T_822; // @[Lookup.scala 33:37]
  wire  _T_823; // @[Lookup.scala 33:37]
  wire  _T_824; // @[Lookup.scala 33:37]
  wire  _T_825; // @[Lookup.scala 33:37]
  wire  _T_826; // @[Lookup.scala 33:37]
  wire  _T_827; // @[Lookup.scala 33:37]
  wire  _T_828; // @[Lookup.scala 33:37]
  wire  _T_829; // @[Lookup.scala 33:37]
  wire  _T_830; // @[Lookup.scala 33:37]
  wire  _T_831; // @[Lookup.scala 33:37]
  wire  _T_832; // @[Lookup.scala 33:37]
  wire  _T_833; // @[Lookup.scala 33:37]
  wire  _T_834; // @[Lookup.scala 33:37]
  wire  _T_835; // @[Lookup.scala 33:37]
  wire  _T_836; // @[Lookup.scala 33:37]
  wire  _T_837; // @[Lookup.scala 33:37]
  wire  _T_838; // @[Lookup.scala 33:37]
  wire  _T_839; // @[Lookup.scala 33:37]
  wire  _T_840; // @[Lookup.scala 33:37]
  wire  _T_841; // @[Lookup.scala 33:37]
  wire [31:0] _T_911; // @[Lookup.scala 33:37]
  wire [31:0] _T_912; // @[Lookup.scala 33:37]
  wire [31:0] _T_913; // @[Lookup.scala 33:37]
  wire [31:0] _T_914; // @[Lookup.scala 33:37]
  wire [31:0] _T_915; // @[Lookup.scala 33:37]
  wire [31:0] _T_916; // @[Lookup.scala 33:37]
  wire [31:0] _T_917; // @[Lookup.scala 33:37]
  wire [31:0] _T_918; // @[Lookup.scala 33:37]
  wire [31:0] _T_919; // @[Lookup.scala 33:37]
  wire [31:0] _T_920; // @[Lookup.scala 33:37]
  wire [31:0] _T_921; // @[Lookup.scala 33:37]
  wire [31:0] _T_922; // @[Lookup.scala 33:37]
  wire [31:0] _T_923; // @[Lookup.scala 33:37]
  wire [31:0] _T_924; // @[Lookup.scala 33:37]
  wire [31:0] _T_925; // @[Lookup.scala 33:37]
  wire [31:0] _T_926; // @[Lookup.scala 33:37]
  wire [31:0] _T_927; // @[Lookup.scala 33:37]
  wire [31:0] _T_928; // @[Lookup.scala 33:37]
  wire [31:0] _T_929; // @[Lookup.scala 33:37]
  wire [31:0] _T_930; // @[Lookup.scala 33:37]
  wire [31:0] _T_931; // @[Lookup.scala 33:37]
  wire [31:0] _T_932; // @[Lookup.scala 33:37]
  wire [31:0] _T_933; // @[Lookup.scala 33:37]
  wire [31:0] _T_934; // @[Lookup.scala 33:37]
  wire [31:0] _T_935; // @[Lookup.scala 33:37]
  wire [31:0] _T_936; // @[Lookup.scala 33:37]
  wire [31:0] _T_937; // @[Lookup.scala 33:37]
  wire [31:0] _T_938; // @[Lookup.scala 33:37]
  wire [31:0] _T_939; // @[Lookup.scala 33:37]
  wire [31:0] _T_940; // @[Lookup.scala 33:37]
  wire [31:0] _T_941; // @[Lookup.scala 33:37]
  wire [31:0] _T_942; // @[Lookup.scala 33:37]
  wire [31:0] _T_943; // @[Lookup.scala 33:37]
  wire [31:0] _T_944; // @[Lookup.scala 33:37]
  wire [31:0] _T_945; // @[Lookup.scala 33:37]
  wire [31:0] _T_946; // @[Lookup.scala 33:37]
  wire [31:0] _T_947; // @[Lookup.scala 33:37]
  wire [31:0] _T_948; // @[Lookup.scala 33:37]
  wire [31:0] _T_949; // @[Lookup.scala 33:37]
  wire [31:0] _T_950; // @[Lookup.scala 33:37]
  wire [31:0] _T_951; // @[Lookup.scala 33:37]
  wire [31:0] _T_952; // @[Lookup.scala 33:37]
  wire [31:0] _T_953; // @[Lookup.scala 33:37]
  wire [31:0] _T_954; // @[Lookup.scala 33:37]
  wire [31:0] _T_955; // @[Lookup.scala 33:37]
  wire [31:0] _T_956; // @[Lookup.scala 33:37]
  wire [31:0] _T_957; // @[Lookup.scala 33:37]
  wire [31:0] _T_958; // @[Lookup.scala 33:37]
  wire [31:0] _T_959; // @[Lookup.scala 33:37]
  wire [31:0] _T_960; // @[Lookup.scala 33:37]
  wire [31:0] _T_961; // @[Lookup.scala 33:37]
  wire [31:0] _T_962; // @[Lookup.scala 33:37]
  wire [31:0] _T_963; // @[Lookup.scala 33:37]
  wire [31:0] _T_964; // @[Lookup.scala 33:37]
  wire [31:0] _T_965; // @[Lookup.scala 33:37]
  wire [31:0] _T_966; // @[Lookup.scala 33:37]
  wire [31:0] _T_967; // @[Lookup.scala 33:37]
  wire [31:0] _T_968; // @[Lookup.scala 33:37]
  wire [31:0] _T_969; // @[Lookup.scala 33:37]
  wire [31:0] _T_970; // @[Lookup.scala 33:37]
  wire [31:0] _T_971; // @[Lookup.scala 33:37]
  wire [31:0] _T_972; // @[Lookup.scala 33:37]
  wire [31:0] _T_973; // @[Lookup.scala 33:37]
  wire [31:0] _T_974; // @[Lookup.scala 33:37]
  wire [31:0] _T_975; // @[Lookup.scala 33:37]
  wire [31:0] _T_976; // @[Lookup.scala 33:37]
  wire [31:0] _T_977; // @[Lookup.scala 33:37]
  wire [31:0] _T_978; // @[Lookup.scala 33:37]
  wire [31:0] _T_979; // @[Lookup.scala 33:37]
  wire [31:0] _T_1012; // @[Lookup.scala 33:37]
  wire [31:0] _T_1013; // @[Lookup.scala 33:37]
  wire [31:0] _T_1014; // @[Lookup.scala 33:37]
  wire [31:0] _T_1015; // @[Lookup.scala 33:37]
  wire [31:0] _T_1016; // @[Lookup.scala 33:37]
  wire [31:0] _T_1017; // @[Lookup.scala 33:37]
  wire [31:0] _T_1018; // @[Lookup.scala 33:37]
  wire [31:0] _T_1019; // @[Lookup.scala 33:37]
  wire [31:0] _T_1020; // @[Lookup.scala 33:37]
  wire [31:0] _T_1021; // @[Lookup.scala 33:37]
  wire [31:0] _T_1022; // @[Lookup.scala 33:37]
  wire [31:0] _T_1023; // @[Lookup.scala 33:37]
  wire [31:0] _T_1024; // @[Lookup.scala 33:37]
  wire [31:0] _T_1025; // @[Lookup.scala 33:37]
  wire [31:0] _T_1026; // @[Lookup.scala 33:37]
  wire [31:0] _T_1027; // @[Lookup.scala 33:37]
  wire [31:0] _T_1028; // @[Lookup.scala 33:37]
  wire [31:0] _T_1029; // @[Lookup.scala 33:37]
  wire [31:0] _T_1030; // @[Lookup.scala 33:37]
  wire [31:0] _T_1031; // @[Lookup.scala 33:37]
  wire [31:0] _T_1032; // @[Lookup.scala 33:37]
  wire [31:0] _T_1033; // @[Lookup.scala 33:37]
  wire [31:0] _T_1034; // @[Lookup.scala 33:37]
  wire [31:0] _T_1035; // @[Lookup.scala 33:37]
  wire [31:0] _T_1036; // @[Lookup.scala 33:37]
  wire [31:0] _T_1037; // @[Lookup.scala 33:37]
  wire [31:0] _T_1038; // @[Lookup.scala 33:37]
  wire [31:0] _T_1039; // @[Lookup.scala 33:37]
  wire [31:0] _T_1040; // @[Lookup.scala 33:37]
  wire [31:0] _T_1041; // @[Lookup.scala 33:37]
  wire [31:0] _T_1042; // @[Lookup.scala 33:37]
  wire [31:0] _T_1043; // @[Lookup.scala 33:37]
  wire [31:0] _T_1044; // @[Lookup.scala 33:37]
  wire [31:0] _T_1045; // @[Lookup.scala 33:37]
  wire [31:0] _T_1046; // @[Lookup.scala 33:37]
  wire [31:0] _T_1047; // @[Lookup.scala 33:37]
  wire [31:0] _T_1048; // @[Lookup.scala 33:37]
  wire  _T_1081; // @[Lookup.scala 33:37]
  wire  _T_1082; // @[Lookup.scala 33:37]
  wire  _T_1083; // @[Lookup.scala 33:37]
  wire  _T_1084; // @[Lookup.scala 33:37]
  wire  _T_1085; // @[Lookup.scala 33:37]
  wire  _T_1086; // @[Lookup.scala 33:37]
  wire  _T_1087; // @[Lookup.scala 33:37]
  wire  _T_1088; // @[Lookup.scala 33:37]
  wire  _T_1089; // @[Lookup.scala 33:37]
  wire  _T_1090; // @[Lookup.scala 33:37]
  wire  _T_1091; // @[Lookup.scala 33:37]
  wire  _T_1092; // @[Lookup.scala 33:37]
  wire  _T_1093; // @[Lookup.scala 33:37]
  wire  _T_1094; // @[Lookup.scala 33:37]
  wire  _T_1095; // @[Lookup.scala 33:37]
  wire  _T_1096; // @[Lookup.scala 33:37]
  wire  _T_1097; // @[Lookup.scala 33:37]
  wire  _T_1098; // @[Lookup.scala 33:37]
  wire  _T_1099; // @[Lookup.scala 33:37]
  wire  _T_1100; // @[Lookup.scala 33:37]
  wire  _T_1101; // @[Lookup.scala 33:37]
  wire  _T_1102; // @[Lookup.scala 33:37]
  wire  _T_1103; // @[Lookup.scala 33:37]
  wire  _T_1104; // @[Lookup.scala 33:37]
  wire  _T_1105; // @[Lookup.scala 33:37]
  wire  _T_1106; // @[Lookup.scala 33:37]
  wire  _T_1107; // @[Lookup.scala 33:37]
  wire  _T_1108; // @[Lookup.scala 33:37]
  wire  _T_1109; // @[Lookup.scala 33:37]
  wire  _T_1110; // @[Lookup.scala 33:37]
  wire  _T_1111; // @[Lookup.scala 33:37]
  wire  _T_1112; // @[Lookup.scala 33:37]
  wire  _T_1113; // @[Lookup.scala 33:37]
  wire  _T_1114; // @[Lookup.scala 33:37]
  wire  _T_1115; // @[Lookup.scala 33:37]
  wire  _T_1116; // @[Lookup.scala 33:37]
  wire  _T_1117; // @[Lookup.scala 33:37]
  wire  _T_1481; // @[Lookup.scala 33:37]
  wire  _T_1554; // @[Lookup.scala 33:37]
  wire  _T_1613; // @[Lookup.scala 33:37]
  wire  _T_1614; // @[Lookup.scala 33:37]
  wire  _T_1615; // @[Lookup.scala 33:37]
  wire  _T_1616; // @[Lookup.scala 33:37]
  wire  _T_1617; // @[Lookup.scala 33:37]
  wire  _T_1618; // @[Lookup.scala 33:37]
  wire  _T_1619; // @[Lookup.scala 33:37]
  wire  _T_1620; // @[Lookup.scala 33:37]
  wire  _T_1621; // @[Lookup.scala 33:37]
  wire  _T_1622; // @[Lookup.scala 33:37]
  wire  _T_1623; // @[Lookup.scala 33:37]
  wire  _T_1624; // @[Lookup.scala 33:37]
  wire  _T_1625; // @[Lookup.scala 33:37]
  wire  _T_1626; // @[Lookup.scala 33:37]
  wire  _T_1627; // @[Lookup.scala 33:37]
  wire  _T_1628; // @[Lookup.scala 33:37]
  wire  _T_1629; // @[Lookup.scala 33:37]
  wire  _T_1630; // @[Lookup.scala 33:37]
  wire  _T_1631; // @[Lookup.scala 33:37]
  wire  _T_1632; // @[Lookup.scala 33:37]
  wire  _T_1633; // @[Lookup.scala 33:37]
  wire  _T_1634; // @[Lookup.scala 33:37]
  wire  _T_1635; // @[Lookup.scala 33:37]
  wire  _T_1636; // @[Lookup.scala 33:37]
  wire  _T_1637; // @[Lookup.scala 33:37]
  wire  _T_1638; // @[Lookup.scala 33:37]
  wire  _T_1639; // @[Lookup.scala 33:37]
  wire  _T_1640; // @[Lookup.scala 33:37]
  wire  _T_1641; // @[Lookup.scala 33:37]
  wire  _T_1642; // @[Lookup.scala 33:37]
  wire  _T_1643; // @[Lookup.scala 33:37]
  wire  _T_1644; // @[Lookup.scala 33:37]
  wire  _T_1645; // @[Lookup.scala 33:37]
  wire  _T_1646; // @[Lookup.scala 33:37]
  wire  _T_1647; // @[Lookup.scala 33:37]
  wire  _T_1648; // @[Lookup.scala 33:37]
  wire  _T_1649; // @[Lookup.scala 33:37]
  wire  _T_1650; // @[Lookup.scala 33:37]
  wire  _T_1651; // @[Lookup.scala 33:37]
  wire  _T_1652; // @[Lookup.scala 33:37]
  wire  _T_1653; // @[Lookup.scala 33:37]
  wire  _T_1654; // @[Lookup.scala 33:37]
  wire  _T_1655; // @[Lookup.scala 33:37]
  wire  _T_1656; // @[Lookup.scala 33:37]
  wire  _T_1657; // @[Lookup.scala 33:37]
  wire  _T_1658; // @[Lookup.scala 33:37]
  wire  _T_1659; // @[Lookup.scala 33:37]
  wire  _T_1660; // @[Lookup.scala 33:37]
  wire  _T_1661; // @[Lookup.scala 33:37]
  wire  _T_1662; // @[Lookup.scala 33:37]
  wire  _T_1663; // @[Lookup.scala 33:37]
  wire  _T_1664; // @[Lookup.scala 33:37]
  wire  _T_1665; // @[Lookup.scala 33:37]
  wire  _T_1666; // @[Lookup.scala 33:37]
  wire  _T_1667; // @[Lookup.scala 33:37]
  wire  _T_1668; // @[Lookup.scala 33:37]
  wire  _T_1669; // @[Lookup.scala 33:37]
  wire  _T_1681; // @[Lookup.scala 33:37]
  wire  _T_1682; // @[Lookup.scala 33:37]
  wire  _T_1683; // @[Lookup.scala 33:37]
  wire  _T_1684; // @[Lookup.scala 33:37]
  wire  _T_1685; // @[Lookup.scala 33:37]
  wire  _T_1686; // @[Lookup.scala 33:37]
  wire  _T_1687; // @[Lookup.scala 33:37]
  wire  _T_1688; // @[Lookup.scala 33:37]
  wire  _T_1689; // @[Lookup.scala 33:37]
  wire  _T_1690; // @[Lookup.scala 33:37]
  wire  _T_1691; // @[Lookup.scala 33:37]
  wire  _T_1692; // @[Lookup.scala 33:37]
  wire  _T_1693; // @[Lookup.scala 33:37]
  wire  _T_1694; // @[Lookup.scala 33:37]
  wire  _T_1695; // @[Lookup.scala 33:37]
  wire  _T_1696; // @[Lookup.scala 33:37]
  wire  _T_1697; // @[Lookup.scala 33:37]
  wire  _T_1698; // @[Lookup.scala 33:37]
  wire  _T_1699; // @[Lookup.scala 33:37]
  wire  _T_1700; // @[Lookup.scala 33:37]
  wire  _T_1701; // @[Lookup.scala 33:37]
  wire  _T_1702; // @[Lookup.scala 33:37]
  wire  _T_1703; // @[Lookup.scala 33:37]
  wire  _T_1704; // @[Lookup.scala 33:37]
  wire  _T_1705; // @[Lookup.scala 33:37]
  wire  _T_1706; // @[Lookup.scala 33:37]
  wire  _T_1707; // @[Lookup.scala 33:37]
  wire  _T_1708; // @[Lookup.scala 33:37]
  wire  _T_1709; // @[Lookup.scala 33:37]
  wire  _T_1710; // @[Lookup.scala 33:37]
  wire  _T_1711; // @[Lookup.scala 33:37]
  wire  _T_1712; // @[Lookup.scala 33:37]
  wire  _T_1713; // @[Lookup.scala 33:37]
  wire  _T_1714; // @[Lookup.scala 33:37]
  wire  _T_1715; // @[Lookup.scala 33:37]
  wire  _T_1716; // @[Lookup.scala 33:37]
  wire  _T_1717; // @[Lookup.scala 33:37]
  wire  _T_1718; // @[Lookup.scala 33:37]
  wire  _T_1719; // @[Lookup.scala 33:37]
  wire  _T_1720; // @[Lookup.scala 33:37]
  wire  _T_1721; // @[Lookup.scala 33:37]
  wire  _T_1722; // @[Lookup.scala 33:37]
  wire  _T_1723; // @[Lookup.scala 33:37]
  wire  _T_1724; // @[Lookup.scala 33:37]
  wire  _T_1725; // @[Lookup.scala 33:37]
  wire  _T_1726; // @[Lookup.scala 33:37]
  wire  _T_1727; // @[Lookup.scala 33:37]
  wire  _T_1728; // @[Lookup.scala 33:37]
  wire  _T_1729; // @[Lookup.scala 33:37]
  wire  _T_1730; // @[Lookup.scala 33:37]
  wire  _T_1731; // @[Lookup.scala 33:37]
  wire  _T_1732; // @[Lookup.scala 33:37]
  wire  _T_1733; // @[Lookup.scala 33:37]
  wire  _T_1734; // @[Lookup.scala 33:37]
  wire  _T_1735; // @[Lookup.scala 33:37]
  wire  _T_1736; // @[Lookup.scala 33:37]
  wire  _T_1737; // @[Lookup.scala 33:37]
  wire  _T_1738; // @[Lookup.scala 33:37]
  wire  _T_1742; // @[IDecode.scala 1016:40]
  wire  _T_1745; // @[IDecode.scala 1018:40]
  wire  _T_1747; // @[IDecode.scala 1018:71]
  wire  _T_1748; // @[IDecode.scala 1018:112]
  wire  _T_1749; // @[IDecode.scala 1018:98]
  wire  _T_1752; // @[IDecode.scala 1021:40]
  wire  _T_1754; // @[IDecode.scala 1021:67]
  wire  _T_1757; // @[IDecode.scala 1023:40]
  wire  _T_1758; // @[IDecode.scala 1023:83]
  wire  _T_1759; // @[IDecode.scala 1023:68]
  wire [31:0] _GEN_93; // @[IDecode.scala 1027:41]
  wire [31:0] _GEN_94; // @[IDecode.scala 1025:40]
  wire [31:0] _GEN_95; // @[IDecode.scala 1023:102]
  wire [31:0] _GEN_96; // @[IDecode.scala 1021:100]
  wire [31:0] _GEN_98; // @[IDecode.scala 1018:131]
  wire [31:0] _GEN_99; // @[IDecode.scala 1016:76]
  wire  _T_1764; // @[IDecode.scala 1037:58]
  wire  _T_1765; // @[IDecode.scala 1037:40]
  wire  _T_1768; // @[IDecode.scala 1039:40]
  wire  _T_1770; // @[IDecode.scala 1039:71]
  wire  _T_1771; // @[IDecode.scala 1039:112]
  wire  _T_1772; // @[IDecode.scala 1039:98]
  wire  _T_1775; // @[IDecode.scala 1042:40]
  wire  _T_1777; // @[IDecode.scala 1042:67]
  wire  _T_1780; // @[IDecode.scala 1044:40]
  wire  _T_1781; // @[IDecode.scala 1044:83]
  wire  _T_1782; // @[IDecode.scala 1044:68]
  wire [31:0] _GEN_103; // @[IDecode.scala 1048:41]
  wire [31:0] _GEN_104; // @[IDecode.scala 1046:40]
  wire [31:0] _GEN_105; // @[IDecode.scala 1044:102]
  wire [31:0] _GEN_106; // @[IDecode.scala 1042:100]
  wire [31:0] _GEN_108; // @[IDecode.scala 1039:131]
  wire [31:0] _GEN_109; // @[IDecode.scala 1037:76]
  assign _T_12 = io_inst_i[31] ? 20'hfffff : 20'h0; // @[Bitwise.scala 71:12]
  assign _T_19 = {_T_12,io_inst_i[31:25]}; // @[Cat.scala 29:58]
  assign _T_27 = io_inst_i[31] ? 19'h7ffff : 19'h0; // @[Bitwise.scala 71:12]
  assign _T_35 = {_T_27,io_inst_i[31],io_inst_i[7],io_inst_i[30:25],io_inst_i[11:8]}; // @[Cat.scala 29:58]
  assign _T_39 = io_inst_i[31] ? 11'h7ff : 11'h0; // @[Bitwise.scala 71:12]
  assign _T_47 = {_T_39,io_inst_i[31],io_inst_i[19:12],io_inst_i[20],io_inst_i[30:21]}; // @[Cat.scala 29:58]
  assign _T_54 = ~io_ex_csr_reg_we_i & ~io_mem_csr_reg_we_i; // @[IDecode.scala 236:44]
  assign _T_56 = _T_54 & ~io_wb_csr_reg_we_i; // @[IDecode.scala 236:89]
  assign _T_59 = io_ex_not_stall_i | io_mem_not_stall_i; // @[IDecode.scala 239:94]
  assign _T_61 = stallreq_for_reg1_loadrelate | stallreq_for_reg2_loadrelate; // @[IDecode.scala 241:46]
  assign _T_62 = _T_61 | stallreq_for_csr_write_relate; // @[IDecode.scala 241:77]
  assign _T_64 = io_ex_aluop_i == 8'he0; // @[IDecode.scala 244:20]
  assign _T_65 = io_ex_aluop_i == 8'he4; // @[IDecode.scala 244:55]
  assign _T_66 = _T_64 | _T_65; // @[IDecode.scala 244:37]
  assign _T_67 = io_ex_aluop_i == 8'he1; // @[IDecode.scala 244:91]
  assign _T_68 = _T_66 | _T_67; // @[IDecode.scala 244:73]
  assign _T_69 = io_ex_aluop_i == 8'he5; // @[IDecode.scala 245:20]
  assign _T_70 = _T_68 | _T_69; // @[IDecode.scala 244:108]
  assign _T_71 = io_ex_aluop_i == 8'he3; // @[IDecode.scala 245:56]
  assign _T_72 = _T_70 | _T_71; // @[IDecode.scala 245:38]
  assign _T_73 = io_ex_aluop_i == 8'hf0; // @[IDecode.scala 245:91]
  assign _T_74 = _T_72 | _T_73; // @[IDecode.scala 245:73]
  assign _T_75 = io_ex_aluop_i == 8'hf8; // @[IDecode.scala 246:20]
  assign _T_76 = _T_74 | _T_75; // @[IDecode.scala 245:108]
  assign _T_77 = io_ex_aluop_i == 8'h41; // @[IDecode.scala 246:55]
  assign _T_78 = _T_76 | _T_77; // @[IDecode.scala 246:37]
  assign _T_79 = io_ex_aluop_i == 8'h40; // @[IDecode.scala 246:97]
  assign _T_80 = _T_78 | _T_79; // @[IDecode.scala 246:79]
  assign _T_81 = io_ex_aluop_i == 8'h44; // @[IDecode.scala 247:20]
  assign _T_82 = _T_80 | _T_81; // @[IDecode.scala 246:120]
  assign _T_83 = io_ex_aluop_i == 8'h4c; // @[IDecode.scala 247:61]
  assign _T_84 = _T_82 | _T_83; // @[IDecode.scala 247:43]
  assign _T_85 = io_ex_aluop_i == 8'h48; // @[IDecode.scala 247:102]
  assign _T_86 = _T_84 | _T_85; // @[IDecode.scala 247:84]
  assign _T_87 = io_ex_aluop_i == 8'h70; // @[IDecode.scala 248:20]
  assign _T_88 = _T_86 | _T_87; // @[IDecode.scala 247:124]
  assign _T_89 = io_ex_aluop_i == 8'h54; // @[IDecode.scala 248:61]
  assign _T_90 = _T_88 | _T_89; // @[IDecode.scala 248:43]
  assign _T_91 = io_ex_aluop_i == 8'h79; // @[IDecode.scala 248:102]
  assign _T_92 = _T_90 | _T_91; // @[IDecode.scala 248:84]
  assign _T_93 = io_ex_aluop_i == 8'h5c; // @[IDecode.scala 249:20]
  assign _T_130 = instvalid | io_csr_protect_i; // @[IDecode.scala 265:56]
  assign _T_131 = 2'h0 == io_prv_i; // @[Conditional.scala 37:30]
  assign _T_132 = 2'h1 == io_prv_i; // @[Conditional.scala 37:30]
  assign _T_133 = 2'h3 == io_prv_i; // @[Conditional.scala 37:30]
  assign _GEN_0 = _T_133 ? excepttype_is_syscall : io_excepttype_i[11]; // @[Conditional.scala 39:67]
  assign _GEN_1 = _T_132 ? excepttype_is_syscall : io_excepttype_i[9]; // @[Conditional.scala 39:67]
  assign _GEN_2 = _T_132 ? io_excepttype_i[11] : _GEN_0; // @[Conditional.scala 39:67]
  assign _GEN_3 = _T_131 ? excepttype_is_syscall : io_excepttype_i[8]; // @[Conditional.scala 40:58]
  assign _GEN_4 = _T_131 ? io_excepttype_i[9] : _GEN_1; // @[Conditional.scala 40:58]
  assign _GEN_5 = _T_131 ? io_excepttype_i[11] : _GEN_2; // @[Conditional.scala 40:58]
  assign _GEN_8 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[1]; // @[IDecode.scala 259:52]
  assign excepttype_b_1 = io_rst_n ? _GEN_8 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_7 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[0]; // @[IDecode.scala 259:52]
  assign excepttype_b_0 = io_rst_n ? _GEN_7 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_10 = io_is_in_delayslot_i ? 1'h0 : excepttype_is_break; // @[IDecode.scala 259:52]
  assign excepttype_b_3 = io_rst_n ? _GEN_10 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_9 = io_is_in_delayslot_i ? 1'h0 : _T_130; // @[IDecode.scala 259:52]
  assign excepttype_b_2 = io_rst_n ? _GEN_9 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_12 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[5]; // @[IDecode.scala 259:52]
  assign excepttype_b_5 = io_rst_n ? _GEN_12 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_11 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[4]; // @[IDecode.scala 259:52]
  assign excepttype_b_4 = io_rst_n ? _GEN_11 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_14 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[7]; // @[IDecode.scala 259:52]
  assign excepttype_b_7 = io_rst_n ? _GEN_14 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_13 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[6]; // @[IDecode.scala 259:52]
  assign excepttype_b_6 = io_rst_n ? _GEN_13 : 1'h0; // @[IDecode.scala 256:32]
  assign _T_140 = {excepttype_b_7,excepttype_b_6,excepttype_b_5,excepttype_b_4,excepttype_b_3,excepttype_b_2,excepttype_b_1,excepttype_b_0}; // @[IDecode.scala 278:35]
  assign _GEN_16 = io_is_in_delayslot_i ? 1'h0 : _GEN_4; // @[IDecode.scala 259:52]
  assign excepttype_b_9 = io_rst_n ? _GEN_16 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_15 = io_is_in_delayslot_i ? 1'h0 : _GEN_3; // @[IDecode.scala 259:52]
  assign excepttype_b_8 = io_rst_n ? _GEN_15 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_18 = io_is_in_delayslot_i ? 1'h0 : _GEN_5; // @[IDecode.scala 259:52]
  assign excepttype_b_11 = io_rst_n ? _GEN_18 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_17 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[10]; // @[IDecode.scala 259:52]
  assign excepttype_b_10 = io_rst_n ? _GEN_17 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_20 = io_is_in_delayslot_i ? 1'h0 : excepttype_is_sret; // @[IDecode.scala 259:52]
  assign excepttype_b_13 = io_rst_n ? _GEN_20 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_19 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[12]; // @[IDecode.scala 259:52]
  assign excepttype_b_12 = io_rst_n ? _GEN_19 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_22 = io_is_in_delayslot_i ? 1'h0 : excepttype_is_mret; // @[IDecode.scala 259:52]
  assign excepttype_b_15 = io_rst_n ? _GEN_22 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_21 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[14]; // @[IDecode.scala 259:52]
  assign excepttype_b_14 = io_rst_n ? _GEN_21 : 1'h0; // @[IDecode.scala 256:32]
  assign _T_148 = {excepttype_b_15,excepttype_b_14,excepttype_b_13,excepttype_b_12,excepttype_b_11,excepttype_b_10,excepttype_b_9,excepttype_b_8,_T_140}; // @[IDecode.scala 278:35]
  assign _GEN_24 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[17]; // @[IDecode.scala 259:52]
  assign excepttype_b_17 = io_rst_n ? _GEN_24 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_23 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[16]; // @[IDecode.scala 259:52]
  assign excepttype_b_16 = io_rst_n ? _GEN_23 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_26 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[19]; // @[IDecode.scala 259:52]
  assign excepttype_b_19 = io_rst_n ? _GEN_26 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_25 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[18]; // @[IDecode.scala 259:52]
  assign excepttype_b_18 = io_rst_n ? _GEN_25 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_28 = io_is_in_delayslot_i ? 1'h0 : excepttype_is_fence_i; // @[IDecode.scala 259:52]
  assign excepttype_b_21 = io_rst_n ? _GEN_28 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_27 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[20]; // @[IDecode.scala 259:52]
  assign excepttype_b_20 = io_rst_n ? _GEN_27 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_30 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[23]; // @[IDecode.scala 259:52]
  assign excepttype_b_23 = io_rst_n ? _GEN_30 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_29 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[22]; // @[IDecode.scala 259:52]
  assign excepttype_b_22 = io_rst_n ? _GEN_29 : 1'h0; // @[IDecode.scala 256:32]
  assign _T_155 = {excepttype_b_23,excepttype_b_22,excepttype_b_21,excepttype_b_20,excepttype_b_19,excepttype_b_18,excepttype_b_17,excepttype_b_16}; // @[IDecode.scala 278:35]
  assign _GEN_32 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[25]; // @[IDecode.scala 259:52]
  assign excepttype_b_25 = io_rst_n ? _GEN_32 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_31 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[24]; // @[IDecode.scala 259:52]
  assign excepttype_b_24 = io_rst_n ? _GEN_31 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_34 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[27]; // @[IDecode.scala 259:52]
  assign excepttype_b_27 = io_rst_n ? _GEN_34 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_33 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[26]; // @[IDecode.scala 259:52]
  assign excepttype_b_26 = io_rst_n ? _GEN_33 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_36 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[29]; // @[IDecode.scala 259:52]
  assign excepttype_b_29 = io_rst_n ? _GEN_36 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_35 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[28]; // @[IDecode.scala 259:52]
  assign excepttype_b_28 = io_rst_n ? _GEN_35 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_38 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[31]; // @[IDecode.scala 259:52]
  assign excepttype_b_31 = io_rst_n ? _GEN_38 : 1'h0; // @[IDecode.scala 256:32]
  assign _GEN_37 = io_is_in_delayslot_i ? 1'h0 : io_excepttype_i[30]; // @[IDecode.scala 259:52]
  assign excepttype_b_30 = io_rst_n ? _GEN_37 : 1'h0; // @[IDecode.scala 256:32]
  assign _T_164 = {excepttype_b_31,excepttype_b_30,excepttype_b_29,excepttype_b_28,excepttype_b_27,excepttype_b_26,excepttype_b_25,excepttype_b_24,_T_155,_T_148}; // @[IDecode.scala 278:35]
  assign _GEN_6 = io_is_in_delayslot_i ? 1'h0 : io_not_stall_i; // @[IDecode.scala 259:52]
  assign _GEN_39 = io_is_in_delayslot_i ? 32'h0 : _T_164; // @[IDecode.scala 259:52]
  assign _T_167 = ~io_rst_n | io_is_in_delayslot_i; // @[IDecode.scala 285:32]
  assign _T_168 = io_excepttype_i != 32'h0; // @[IDecode.scala 285:93]
  assign _T_170 = _T_167 | _T_168; // @[IDecode.scala 285:74]
  assign _T_172 = imm_u_type + io_pc_i; // @[IDecode.scala 444:19]
  assign _T_174 = io_pc_i + imm_uj_type; // @[IDecode.scala 620:16]
  assign _T_176 = io_reg1_o + imm_i_type; // @[IDecode.scala 629:32]
  assign _T_178 = {1'h0,_T_176[30:0]}; // @[Cat.scala 29:58]
  assign _T_179 = io_reg1_o == io_reg2_o; // @[IDecode.scala 639:23]
  assign _T_181 = io_pc_i + imm_sb_type; // @[IDecode.scala 639:46]
  assign _T_182 = _T_179 ? _T_181 : 32'h0; // @[IDecode.scala 639:12]
  assign _T_187 = io_reg1_o != io_reg2_o; // @[IDecode.scala 648:23]
  assign _T_190 = _T_187 ? _T_181 : 32'h0; // @[IDecode.scala 648:12]
  assign _T_197 = $signed(io_reg1_o) < $signed(io_reg2_o); // @[IDecode.scala 657:30]
  assign _T_200 = _T_197 ? _T_181 : 32'h0; // @[IDecode.scala 657:12]
  assign _T_209 = io_reg1_o < io_reg2_o; // @[IDecode.scala 666:23]
  assign _T_212 = _T_209 ? _T_181 : 32'h0; // @[IDecode.scala 666:12]
  assign _T_219 = $signed(io_reg1_o) >= $signed(io_reg2_o); // @[IDecode.scala 675:30]
  assign _T_222 = _T_219 ? _T_181 : 32'h0; // @[IDecode.scala 675:12]
  assign _T_231 = io_reg1_o >= io_reg2_o; // @[IDecode.scala 684:23]
  assign _T_234 = _T_231 ? _T_181 : 32'h0; // @[IDecode.scala 684:12]
  assign _T_240 = imm_i_type + io_reg1_o; // @[IDecode.scala 693:21]
  assign _T_250 = imm_s_type + io_reg1_o; // @[IDecode.scala 739:21]
  assign _T_255 = io_reg1_addr_o == 5'h0; // @[IDecode.scala 764:60]
  assign _T_256 = io_wd_o == 5'h0; // @[IDecode.scala 764:89]
  assign _T_257 = _T_255 & _T_256; // @[IDecode.scala 764:78]
  assign _T_259 = io_inst_i[31:28] == 4'h0; // @[IDecode.scala 764:127]
  assign _T_260 = _T_257 & _T_259; // @[IDecode.scala 764:107]
  assign _T_265 = imm_i_type == 32'h0; // @[IDecode.scala 773:121]
  assign _T_266 = _T_257 & _T_265; // @[IDecode.scala 773:107]
  assign _T_274 = io_prv_i >= 2'h3; // @[IDecode.scala 810:54]
  assign _T_278 = io_wd_o != 5'h0; // @[IDecode.scala 835:21]
  assign _T_280 = io_reg1_addr_o != 5'h0; // @[IDecode.scala 844:42]
  assign _T_290 = io_inst_i & 32'h707f; // @[Lookup.scala 31:38]
  assign _T_291 = 32'h13 == _T_290; // @[Lookup.scala 31:38]
  assign _T_293 = 32'h2013 == _T_290; // @[Lookup.scala 31:38]
  assign _T_295 = 32'h3013 == _T_290; // @[Lookup.scala 31:38]
  assign _T_297 = 32'h7013 == _T_290; // @[Lookup.scala 31:38]
  assign _T_299 = 32'h6013 == _T_290; // @[Lookup.scala 31:38]
  assign _T_301 = 32'h4013 == _T_290; // @[Lookup.scala 31:38]
  assign _T_302 = io_inst_i & 32'hfc00707f; // @[Lookup.scala 31:38]
  assign _T_303 = 32'h1013 == _T_302; // @[Lookup.scala 31:38]
  assign _T_305 = 32'h5013 == _T_302; // @[Lookup.scala 31:38]
  assign _T_307 = 32'h40005013 == _T_302; // @[Lookup.scala 31:38]
  assign _T_308 = io_inst_i & 32'h7f; // @[Lookup.scala 31:38]
  assign _T_309 = 32'h37 == _T_308; // @[Lookup.scala 31:38]
  assign _T_311 = 32'h17 == _T_308; // @[Lookup.scala 31:38]
  assign _T_312 = io_inst_i & 32'hfe00707f; // @[Lookup.scala 31:38]
  assign _T_313 = 32'h33 == _T_312; // @[Lookup.scala 31:38]
  assign _T_315 = 32'h40000033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_317 = 32'h2000033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_319 = 32'h1033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_321 = 32'h2001033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_323 = 32'h2033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_325 = 32'h2002033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_327 = 32'h3033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_329 = 32'h2003033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_331 = 32'h4033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_333 = 32'h2004033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_335 = 32'h5033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_337 = 32'h40005033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_339 = 32'h2005033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_341 = 32'h6033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_343 = 32'h2006033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_345 = 32'h7033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_347 = 32'h2007033 == _T_312; // @[Lookup.scala 31:38]
  assign _T_349 = 32'h6f == _T_308; // @[Lookup.scala 31:38]
  assign _T_351 = 32'h67 == _T_290; // @[Lookup.scala 31:38]
  assign _T_353 = 32'h63 == _T_290; // @[Lookup.scala 31:38]
  assign _T_355 = 32'h1063 == _T_290; // @[Lookup.scala 31:38]
  assign _T_357 = 32'h4063 == _T_290; // @[Lookup.scala 31:38]
  assign _T_359 = 32'h6063 == _T_290; // @[Lookup.scala 31:38]
  assign _T_361 = 32'h5063 == _T_290; // @[Lookup.scala 31:38]
  assign _T_363 = 32'h7063 == _T_290; // @[Lookup.scala 31:38]
  assign _T_365 = 32'h3 == _T_290; // @[Lookup.scala 31:38]
  assign _T_367 = 32'h1003 == _T_290; // @[Lookup.scala 31:38]
  assign _T_369 = 32'h2003 == _T_290; // @[Lookup.scala 31:38]
  assign _T_371 = 32'h4003 == _T_290; // @[Lookup.scala 31:38]
  assign _T_373 = 32'h5003 == _T_290; // @[Lookup.scala 31:38]
  assign _T_375 = 32'h23 == _T_290; // @[Lookup.scala 31:38]
  assign _T_377 = 32'h1023 == _T_290; // @[Lookup.scala 31:38]
  assign _T_379 = 32'h2023 == _T_290; // @[Lookup.scala 31:38]
  assign _T_381 = 32'hf == _T_290; // @[Lookup.scala 31:38]
  assign _T_383 = 32'h100f == io_inst_i; // @[Lookup.scala 31:38]
  assign _T_385 = 32'h73 == io_inst_i; // @[Lookup.scala 31:38]
  assign _T_387 = 32'h100073 == io_inst_i; // @[Lookup.scala 31:38]
  assign _T_389 = 32'h10200073 == io_inst_i; // @[Lookup.scala 31:38]
  assign _T_391 = 32'h30200073 == io_inst_i; // @[Lookup.scala 31:38]
  assign _T_393 = 32'h10500073 == io_inst_i; // @[Lookup.scala 31:38]
  assign _T_395 = 32'h1073 == _T_290; // @[Lookup.scala 31:38]
  assign _T_397 = 32'h2073 == _T_290; // @[Lookup.scala 31:38]
  assign _T_399 = 32'h3073 == _T_290; // @[Lookup.scala 31:38]
  assign _T_401 = 32'h5073 == _T_290; // @[Lookup.scala 31:38]
  assign _T_403 = 32'h6073 == _T_290; // @[Lookup.scala 31:38]
  assign _T_405 = 32'h7073 == _T_290; // @[Lookup.scala 31:38]
  assign _T_406 = io_inst_i & 32'hf9f0707f; // @[Lookup.scala 31:38]
  assign _T_407 = 32'h1000202f == _T_406; // @[Lookup.scala 31:38]
  assign _T_408 = io_inst_i & 32'hf800707f; // @[Lookup.scala 31:38]
  assign _T_409 = 32'h1800202f == _T_408; // @[Lookup.scala 31:38]
  assign _T_411 = 32'h800202f == _T_408; // @[Lookup.scala 31:38]
  assign _T_413 = 32'h202f == _T_408; // @[Lookup.scala 31:38]
  assign _T_415 = 32'h2000202f == _T_408; // @[Lookup.scala 31:38]
  assign _T_417 = 32'h6000202f == _T_408; // @[Lookup.scala 31:38]
  assign _T_419 = 32'h4000202f == _T_408; // @[Lookup.scala 31:38]
  assign _T_421 = 32'h8000202f == _T_408; // @[Lookup.scala 31:38]
  assign _T_423 = 32'ha000202f == _T_408; // @[Lookup.scala 31:38]
  assign _T_425 = 32'hc000202f == _T_408; // @[Lookup.scala 31:38]
  assign _T_427 = 32'he000202f == _T_408; // @[Lookup.scala 31:38]
  assign _T_428 = _T_427 ? 8'h5c : 8'h0; // @[Lookup.scala 33:37]
  assign _T_429 = _T_425 ? 8'h79 : _T_428; // @[Lookup.scala 33:37]
  assign _T_430 = _T_423 ? 8'h54 : _T_429; // @[Lookup.scala 33:37]
  assign _T_431 = _T_421 ? 8'h70 : _T_430; // @[Lookup.scala 33:37]
  assign _T_432 = _T_419 ? 8'h48 : _T_431; // @[Lookup.scala 33:37]
  assign _T_433 = _T_417 ? 8'h4c : _T_432; // @[Lookup.scala 33:37]
  assign _T_434 = _T_415 ? 8'h44 : _T_433; // @[Lookup.scala 33:37]
  assign _T_435 = _T_413 ? 8'h40 : _T_434; // @[Lookup.scala 33:37]
  assign _T_436 = _T_411 ? 8'h41 : _T_435; // @[Lookup.scala 33:37]
  assign _T_437 = _T_409 ? 8'hf8 : _T_436; // @[Lookup.scala 33:37]
  assign _T_438 = _T_407 ? 8'hf0 : _T_437; // @[Lookup.scala 33:37]
  assign _T_439 = _T_405 ? 8'h5a : _T_438; // @[Lookup.scala 33:37]
  assign _T_440 = _T_403 ? 8'h59 : _T_439; // @[Lookup.scala 33:37]
  assign _T_441 = _T_401 ? 8'h58 : _T_440; // @[Lookup.scala 33:37]
  assign _T_442 = _T_399 ? 8'h5a : _T_441; // @[Lookup.scala 33:37]
  assign _T_443 = _T_397 ? 8'h59 : _T_442; // @[Lookup.scala 33:37]
  assign _T_444 = _T_395 ? 8'h58 : _T_443; // @[Lookup.scala 33:37]
  assign _T_445 = _T_393 ? 8'h0 : _T_444; // @[Lookup.scala 33:37]
  assign _T_446 = _T_391 ? 8'h0 : _T_445; // @[Lookup.scala 33:37]
  assign _T_447 = _T_389 ? 8'h0 : _T_446; // @[Lookup.scala 33:37]
  assign _T_448 = _T_387 ? 8'h0 : _T_447; // @[Lookup.scala 33:37]
  assign _T_449 = _T_385 ? 8'h0 : _T_448; // @[Lookup.scala 33:37]
  assign _T_450 = _T_383 ? 8'h0 : _T_449; // @[Lookup.scala 33:37]
  assign _T_451 = _T_381 ? 8'h0 : _T_450; // @[Lookup.scala 33:37]
  assign _T_452 = _T_379 ? 8'heb : _T_451; // @[Lookup.scala 33:37]
  assign _T_453 = _T_377 ? 8'he9 : _T_452; // @[Lookup.scala 33:37]
  assign _T_454 = _T_375 ? 8'he8 : _T_453; // @[Lookup.scala 33:37]
  assign _T_455 = _T_373 ? 8'he5 : _T_454; // @[Lookup.scala 33:37]
  assign _T_456 = _T_371 ? 8'he4 : _T_455; // @[Lookup.scala 33:37]
  assign _T_457 = _T_369 ? 8'he3 : _T_456; // @[Lookup.scala 33:37]
  assign _T_458 = _T_367 ? 8'he1 : _T_457; // @[Lookup.scala 33:37]
  assign _T_459 = _T_365 ? 8'he0 : _T_458; // @[Lookup.scala 33:37]
  assign _T_460 = _T_363 ? 8'h0 : _T_459; // @[Lookup.scala 33:37]
  assign _T_461 = _T_361 ? 8'h0 : _T_460; // @[Lookup.scala 33:37]
  assign _T_462 = _T_359 ? 8'h0 : _T_461; // @[Lookup.scala 33:37]
  assign _T_463 = _T_357 ? 8'h0 : _T_462; // @[Lookup.scala 33:37]
  assign _T_464 = _T_355 ? 8'h0 : _T_463; // @[Lookup.scala 33:37]
  assign _T_465 = _T_353 ? 8'h0 : _T_464; // @[Lookup.scala 33:37]
  assign _T_466 = _T_351 ? 8'h50 : _T_465; // @[Lookup.scala 33:37]
  assign _T_467 = _T_349 ? 8'h50 : _T_466; // @[Lookup.scala 33:37]
  assign _T_468 = _T_347 ? 8'haa : _T_467; // @[Lookup.scala 33:37]
  assign _T_469 = _T_345 ? 8'h24 : _T_468; // @[Lookup.scala 33:37]
  assign _T_470 = _T_343 ? 8'ha8 : _T_469; // @[Lookup.scala 33:37]
  assign _T_471 = _T_341 ? 8'h25 : _T_470; // @[Lookup.scala 33:37]
  assign _T_472 = _T_339 ? 8'h1b : _T_471; // @[Lookup.scala 33:37]
  assign _T_473 = _T_337 ? 8'h3 : _T_472; // @[Lookup.scala 33:37]
  assign _T_474 = _T_335 ? 8'h2 : _T_473; // @[Lookup.scala 33:37]
  assign _T_475 = _T_333 ? 8'h1a : _T_474; // @[Lookup.scala 33:37]
  assign _T_476 = _T_331 ? 8'h26 : _T_475; // @[Lookup.scala 33:37]
  assign _T_477 = _T_329 ? 8'ha6 : _T_476; // @[Lookup.scala 33:37]
  assign _T_478 = _T_327 ? 8'h2b : _T_477; // @[Lookup.scala 33:37]
  assign _T_479 = _T_325 ? 8'ha9 : _T_478; // @[Lookup.scala 33:37]
  assign _T_480 = _T_323 ? 8'h2a : _T_479; // @[Lookup.scala 33:37]
  assign _T_481 = _T_321 ? 8'h19 : _T_480; // @[Lookup.scala 33:37]
  assign _T_482 = _T_319 ? 8'h7c : _T_481; // @[Lookup.scala 33:37]
  assign _T_483 = _T_317 ? 8'h18 : _T_482; // @[Lookup.scala 33:37]
  assign _T_484 = _T_315 ? 8'h22 : _T_483; // @[Lookup.scala 33:37]
  assign _T_485 = _T_313 ? 8'h20 : _T_484; // @[Lookup.scala 33:37]
  assign _T_486 = _T_311 ? 8'h25 : _T_485; // @[Lookup.scala 33:37]
  assign _T_487 = _T_309 ? 8'h25 : _T_486; // @[Lookup.scala 33:37]
  assign _T_488 = _T_307 ? 8'h3 : _T_487; // @[Lookup.scala 33:37]
  assign _T_489 = _T_305 ? 8'h2 : _T_488; // @[Lookup.scala 33:37]
  assign _T_490 = _T_303 ? 8'h7c : _T_489; // @[Lookup.scala 33:37]
  assign _T_491 = _T_301 ? 8'h26 : _T_490; // @[Lookup.scala 33:37]
  assign _T_492 = _T_299 ? 8'h25 : _T_491; // @[Lookup.scala 33:37]
  assign _T_493 = _T_297 ? 8'h24 : _T_492; // @[Lookup.scala 33:37]
  assign _T_494 = _T_295 ? 8'h2b : _T_493; // @[Lookup.scala 33:37]
  assign _T_495 = _T_293 ? 8'h2a : _T_494; // @[Lookup.scala 33:37]
  assign _T_496 = _T_291 ? 8'h20 : _T_495; // @[Lookup.scala 33:37]
  assign _T_497 = _T_427 ? 3'h7 : 3'h0; // @[Lookup.scala 33:37]
  assign _T_498 = _T_425 ? 3'h7 : _T_497; // @[Lookup.scala 33:37]
  assign _T_499 = _T_423 ? 3'h7 : _T_498; // @[Lookup.scala 33:37]
  assign _T_500 = _T_421 ? 3'h7 : _T_499; // @[Lookup.scala 33:37]
  assign _T_501 = _T_419 ? 3'h7 : _T_500; // @[Lookup.scala 33:37]
  assign _T_502 = _T_417 ? 3'h7 : _T_501; // @[Lookup.scala 33:37]
  assign _T_503 = _T_415 ? 3'h7 : _T_502; // @[Lookup.scala 33:37]
  assign _T_504 = _T_413 ? 3'h7 : _T_503; // @[Lookup.scala 33:37]
  assign _T_505 = _T_411 ? 3'h7 : _T_504; // @[Lookup.scala 33:37]
  assign _T_506 = _T_409 ? 3'h7 : _T_505; // @[Lookup.scala 33:37]
  assign _T_507 = _T_407 ? 3'h7 : _T_506; // @[Lookup.scala 33:37]
  assign _T_508 = _T_405 ? 3'h3 : _T_507; // @[Lookup.scala 33:37]
  assign _T_509 = _T_403 ? 3'h3 : _T_508; // @[Lookup.scala 33:37]
  assign _T_510 = _T_401 ? 3'h3 : _T_509; // @[Lookup.scala 33:37]
  assign _T_511 = _T_399 ? 3'h3 : _T_510; // @[Lookup.scala 33:37]
  assign _T_512 = _T_397 ? 3'h3 : _T_511; // @[Lookup.scala 33:37]
  assign _T_513 = _T_395 ? 3'h3 : _T_512; // @[Lookup.scala 33:37]
  assign _T_514 = _T_393 ? 3'h0 : _T_513; // @[Lookup.scala 33:37]
  assign _T_515 = _T_391 ? 3'h0 : _T_514; // @[Lookup.scala 33:37]
  assign _T_516 = _T_389 ? 3'h0 : _T_515; // @[Lookup.scala 33:37]
  assign _T_517 = _T_387 ? 3'h0 : _T_516; // @[Lookup.scala 33:37]
  assign _T_518 = _T_385 ? 3'h0 : _T_517; // @[Lookup.scala 33:37]
  assign _T_519 = _T_383 ? 3'h0 : _T_518; // @[Lookup.scala 33:37]
  assign _T_520 = _T_381 ? 3'h0 : _T_519; // @[Lookup.scala 33:37]
  assign _T_521 = _T_379 ? 3'h7 : _T_520; // @[Lookup.scala 33:37]
  assign _T_522 = _T_377 ? 3'h7 : _T_521; // @[Lookup.scala 33:37]
  assign _T_523 = _T_375 ? 3'h7 : _T_522; // @[Lookup.scala 33:37]
  assign _T_524 = _T_373 ? 3'h7 : _T_523; // @[Lookup.scala 33:37]
  assign _T_525 = _T_371 ? 3'h7 : _T_524; // @[Lookup.scala 33:37]
  assign _T_526 = _T_369 ? 3'h7 : _T_525; // @[Lookup.scala 33:37]
  assign _T_527 = _T_367 ? 3'h7 : _T_526; // @[Lookup.scala 33:37]
  assign _T_528 = _T_365 ? 3'h7 : _T_527; // @[Lookup.scala 33:37]
  assign _T_529 = _T_363 ? 3'h0 : _T_528; // @[Lookup.scala 33:37]
  assign _T_530 = _T_361 ? 3'h0 : _T_529; // @[Lookup.scala 33:37]
  assign _T_531 = _T_359 ? 3'h0 : _T_530; // @[Lookup.scala 33:37]
  assign _T_532 = _T_357 ? 3'h0 : _T_531; // @[Lookup.scala 33:37]
  assign _T_533 = _T_355 ? 3'h0 : _T_532; // @[Lookup.scala 33:37]
  assign _T_534 = _T_353 ? 3'h0 : _T_533; // @[Lookup.scala 33:37]
  assign _T_535 = _T_351 ? 3'h6 : _T_534; // @[Lookup.scala 33:37]
  assign _T_536 = _T_349 ? 3'h6 : _T_535; // @[Lookup.scala 33:37]
  assign _T_537 = _T_347 ? 3'h5 : _T_536; // @[Lookup.scala 33:37]
  assign _T_538 = _T_345 ? 3'h1 : _T_537; // @[Lookup.scala 33:37]
  assign _T_539 = _T_343 ? 3'h5 : _T_538; // @[Lookup.scala 33:37]
  assign _T_540 = _T_341 ? 3'h1 : _T_539; // @[Lookup.scala 33:37]
  assign _T_541 = _T_339 ? 3'h5 : _T_540; // @[Lookup.scala 33:37]
  assign _T_542 = _T_337 ? 3'h2 : _T_541; // @[Lookup.scala 33:37]
  assign _T_543 = _T_335 ? 3'h2 : _T_542; // @[Lookup.scala 33:37]
  assign _T_544 = _T_333 ? 3'h5 : _T_543; // @[Lookup.scala 33:37]
  assign _T_545 = _T_331 ? 3'h1 : _T_544; // @[Lookup.scala 33:37]
  assign _T_546 = _T_329 ? 3'h5 : _T_545; // @[Lookup.scala 33:37]
  assign _T_547 = _T_327 ? 3'h4 : _T_546; // @[Lookup.scala 33:37]
  assign _T_548 = _T_325 ? 3'h5 : _T_547; // @[Lookup.scala 33:37]
  assign _T_549 = _T_323 ? 3'h4 : _T_548; // @[Lookup.scala 33:37]
  assign _T_550 = _T_321 ? 3'h5 : _T_549; // @[Lookup.scala 33:37]
  assign _T_551 = _T_319 ? 3'h2 : _T_550; // @[Lookup.scala 33:37]
  assign _T_552 = _T_317 ? 3'h5 : _T_551; // @[Lookup.scala 33:37]
  assign _T_553 = _T_315 ? 3'h4 : _T_552; // @[Lookup.scala 33:37]
  assign _T_554 = _T_313 ? 3'h4 : _T_553; // @[Lookup.scala 33:37]
  assign _T_555 = _T_311 ? 3'h1 : _T_554; // @[Lookup.scala 33:37]
  assign _T_556 = _T_309 ? 3'h1 : _T_555; // @[Lookup.scala 33:37]
  assign _T_557 = _T_307 ? 3'h2 : _T_556; // @[Lookup.scala 33:37]
  assign _T_558 = _T_305 ? 3'h2 : _T_557; // @[Lookup.scala 33:37]
  assign _T_559 = _T_303 ? 3'h2 : _T_558; // @[Lookup.scala 33:37]
  assign _T_560 = _T_301 ? 3'h1 : _T_559; // @[Lookup.scala 33:37]
  assign _T_561 = _T_299 ? 3'h1 : _T_560; // @[Lookup.scala 33:37]
  assign _T_562 = _T_297 ? 3'h1 : _T_561; // @[Lookup.scala 33:37]
  assign _T_563 = _T_295 ? 3'h4 : _T_562; // @[Lookup.scala 33:37]
  assign _T_564 = _T_293 ? 3'h4 : _T_563; // @[Lookup.scala 33:37]
  assign _T_565 = _T_291 ? 3'h4 : _T_564; // @[Lookup.scala 33:37]
  assign _T_636 = _T_425 | _T_427; // @[Lookup.scala 33:37]
  assign _T_637 = _T_423 | _T_636; // @[Lookup.scala 33:37]
  assign _T_638 = _T_421 | _T_637; // @[Lookup.scala 33:37]
  assign _T_639 = _T_419 | _T_638; // @[Lookup.scala 33:37]
  assign _T_640 = _T_417 | _T_639; // @[Lookup.scala 33:37]
  assign _T_641 = _T_415 | _T_640; // @[Lookup.scala 33:37]
  assign _T_642 = _T_413 | _T_641; // @[Lookup.scala 33:37]
  assign _T_643 = _T_411 | _T_642; // @[Lookup.scala 33:37]
  assign _T_644 = _T_409 | _T_643; // @[Lookup.scala 33:37]
  assign _T_645 = _T_407 | _T_644; // @[Lookup.scala 33:37]
  assign _T_646 = _T_405 | _T_645; // @[Lookup.scala 33:37]
  assign _T_647 = _T_403 | _T_646; // @[Lookup.scala 33:37]
  assign _T_648 = _T_401 | _T_647; // @[Lookup.scala 33:37]
  assign _T_649 = _T_399 | _T_648; // @[Lookup.scala 33:37]
  assign _T_650 = _T_397 | _T_649; // @[Lookup.scala 33:37]
  assign _T_651 = _T_395 | _T_650; // @[Lookup.scala 33:37]
  assign _T_652 = _T_393 ? 1'h0 : _T_651; // @[Lookup.scala 33:37]
  assign _T_653 = _T_391 ? 1'h0 : _T_652; // @[Lookup.scala 33:37]
  assign _T_654 = _T_389 ? 1'h0 : _T_653; // @[Lookup.scala 33:37]
  assign _T_655 = _T_387 ? 1'h0 : _T_654; // @[Lookup.scala 33:37]
  assign _T_656 = _T_385 ? 1'h0 : _T_655; // @[Lookup.scala 33:37]
  assign _T_657 = _T_383 ? 1'h0 : _T_656; // @[Lookup.scala 33:37]
  assign _T_658 = _T_381 ? 1'h0 : _T_657; // @[Lookup.scala 33:37]
  assign _T_659 = _T_379 ? 1'h0 : _T_658; // @[Lookup.scala 33:37]
  assign _T_660 = _T_377 ? 1'h0 : _T_659; // @[Lookup.scala 33:37]
  assign _T_661 = _T_375 ? 1'h0 : _T_660; // @[Lookup.scala 33:37]
  assign _T_662 = _T_373 | _T_661; // @[Lookup.scala 33:37]
  assign _T_663 = _T_371 | _T_662; // @[Lookup.scala 33:37]
  assign _T_664 = _T_369 | _T_663; // @[Lookup.scala 33:37]
  assign _T_665 = _T_367 | _T_664; // @[Lookup.scala 33:37]
  assign _T_666 = _T_365 | _T_665; // @[Lookup.scala 33:37]
  assign _T_667 = _T_363 ? 1'h0 : _T_666; // @[Lookup.scala 33:37]
  assign _T_668 = _T_361 ? 1'h0 : _T_667; // @[Lookup.scala 33:37]
  assign _T_669 = _T_359 ? 1'h0 : _T_668; // @[Lookup.scala 33:37]
  assign _T_670 = _T_357 ? 1'h0 : _T_669; // @[Lookup.scala 33:37]
  assign _T_671 = _T_355 ? 1'h0 : _T_670; // @[Lookup.scala 33:37]
  assign _T_672 = _T_353 ? 1'h0 : _T_671; // @[Lookup.scala 33:37]
  assign _T_673 = _T_351 | _T_672; // @[Lookup.scala 33:37]
  assign _T_674 = _T_349 | _T_673; // @[Lookup.scala 33:37]
  assign _T_675 = _T_347 | _T_674; // @[Lookup.scala 33:37]
  assign _T_676 = _T_345 | _T_675; // @[Lookup.scala 33:37]
  assign _T_677 = _T_343 | _T_676; // @[Lookup.scala 33:37]
  assign _T_678 = _T_341 | _T_677; // @[Lookup.scala 33:37]
  assign _T_679 = _T_339 | _T_678; // @[Lookup.scala 33:37]
  assign _T_680 = _T_337 | _T_679; // @[Lookup.scala 33:37]
  assign _T_681 = _T_335 | _T_680; // @[Lookup.scala 33:37]
  assign _T_682 = _T_333 | _T_681; // @[Lookup.scala 33:37]
  assign _T_683 = _T_331 | _T_682; // @[Lookup.scala 33:37]
  assign _T_684 = _T_329 | _T_683; // @[Lookup.scala 33:37]
  assign _T_685 = _T_327 | _T_684; // @[Lookup.scala 33:37]
  assign _T_686 = _T_325 | _T_685; // @[Lookup.scala 33:37]
  assign _T_687 = _T_323 | _T_686; // @[Lookup.scala 33:37]
  assign _T_688 = _T_321 | _T_687; // @[Lookup.scala 33:37]
  assign _T_689 = _T_319 | _T_688; // @[Lookup.scala 33:37]
  assign _T_690 = _T_317 | _T_689; // @[Lookup.scala 33:37]
  assign _T_691 = _T_315 | _T_690; // @[Lookup.scala 33:37]
  assign _T_692 = _T_313 | _T_691; // @[Lookup.scala 33:37]
  assign _T_693 = _T_311 | _T_692; // @[Lookup.scala 33:37]
  assign _T_694 = _T_309 | _T_693; // @[Lookup.scala 33:37]
  assign _T_695 = _T_307 | _T_694; // @[Lookup.scala 33:37]
  assign _T_696 = _T_305 | _T_695; // @[Lookup.scala 33:37]
  assign _T_697 = _T_303 | _T_696; // @[Lookup.scala 33:37]
  assign _T_698 = _T_301 | _T_697; // @[Lookup.scala 33:37]
  assign _T_699 = _T_299 | _T_698; // @[Lookup.scala 33:37]
  assign _T_700 = _T_297 | _T_699; // @[Lookup.scala 33:37]
  assign _T_701 = _T_295 | _T_700; // @[Lookup.scala 33:37]
  assign _T_702 = _T_293 | _T_701; // @[Lookup.scala 33:37]
  assign _T_703 = _T_291 | _T_702; // @[Lookup.scala 33:37]
  assign _T_728 = _T_379 | _T_658; // @[Lookup.scala 33:37]
  assign _T_729 = _T_377 | _T_728; // @[Lookup.scala 33:37]
  assign _T_730 = _T_375 | _T_729; // @[Lookup.scala 33:37]
  assign _T_731 = _T_373 | _T_730; // @[Lookup.scala 33:37]
  assign _T_732 = _T_371 | _T_731; // @[Lookup.scala 33:37]
  assign _T_733 = _T_369 | _T_732; // @[Lookup.scala 33:37]
  assign _T_734 = _T_367 | _T_733; // @[Lookup.scala 33:37]
  assign _T_735 = _T_365 | _T_734; // @[Lookup.scala 33:37]
  assign _T_736 = _T_363 | _T_735; // @[Lookup.scala 33:37]
  assign _T_737 = _T_361 | _T_736; // @[Lookup.scala 33:37]
  assign _T_738 = _T_359 | _T_737; // @[Lookup.scala 33:37]
  assign _T_739 = _T_357 | _T_738; // @[Lookup.scala 33:37]
  assign _T_740 = _T_355 | _T_739; // @[Lookup.scala 33:37]
  assign _T_741 = _T_353 | _T_740; // @[Lookup.scala 33:37]
  assign _T_742 = _T_351 | _T_741; // @[Lookup.scala 33:37]
  assign _T_743 = _T_349 ? 1'h0 : _T_742; // @[Lookup.scala 33:37]
  assign _T_744 = _T_347 | _T_743; // @[Lookup.scala 33:37]
  assign _T_745 = _T_345 | _T_744; // @[Lookup.scala 33:37]
  assign _T_746 = _T_343 | _T_745; // @[Lookup.scala 33:37]
  assign _T_747 = _T_341 | _T_746; // @[Lookup.scala 33:37]
  assign _T_748 = _T_339 | _T_747; // @[Lookup.scala 33:37]
  assign _T_749 = _T_337 | _T_748; // @[Lookup.scala 33:37]
  assign _T_750 = _T_335 | _T_749; // @[Lookup.scala 33:37]
  assign _T_751 = _T_333 | _T_750; // @[Lookup.scala 33:37]
  assign _T_752 = _T_331 | _T_751; // @[Lookup.scala 33:37]
  assign _T_753 = _T_329 | _T_752; // @[Lookup.scala 33:37]
  assign _T_754 = _T_327 | _T_753; // @[Lookup.scala 33:37]
  assign _T_755 = _T_325 | _T_754; // @[Lookup.scala 33:37]
  assign _T_756 = _T_323 | _T_755; // @[Lookup.scala 33:37]
  assign _T_757 = _T_321 | _T_756; // @[Lookup.scala 33:37]
  assign _T_758 = _T_319 | _T_757; // @[Lookup.scala 33:37]
  assign _T_759 = _T_317 | _T_758; // @[Lookup.scala 33:37]
  assign _T_760 = _T_315 | _T_759; // @[Lookup.scala 33:37]
  assign _T_761 = _T_313 | _T_760; // @[Lookup.scala 33:37]
  assign _T_762 = _T_311 ? 1'h0 : _T_761; // @[Lookup.scala 33:37]
  assign _T_763 = _T_309 ? 1'h0 : _T_762; // @[Lookup.scala 33:37]
  assign _T_764 = _T_307 | _T_763; // @[Lookup.scala 33:37]
  assign _T_765 = _T_305 | _T_764; // @[Lookup.scala 33:37]
  assign _T_766 = _T_303 | _T_765; // @[Lookup.scala 33:37]
  assign _T_767 = _T_301 | _T_766; // @[Lookup.scala 33:37]
  assign _T_768 = _T_299 | _T_767; // @[Lookup.scala 33:37]
  assign _T_769 = _T_297 | _T_768; // @[Lookup.scala 33:37]
  assign _T_770 = _T_295 | _T_769; // @[Lookup.scala 33:37]
  assign _T_771 = _T_293 | _T_770; // @[Lookup.scala 33:37]
  assign _T_772 = _T_291 | _T_771; // @[Lookup.scala 33:37]
  assign _T_783 = _T_407 ? 1'h0 : _T_644; // @[Lookup.scala 33:37]
  assign _T_784 = _T_405 ? 1'h0 : _T_783; // @[Lookup.scala 33:37]
  assign _T_785 = _T_403 ? 1'h0 : _T_784; // @[Lookup.scala 33:37]
  assign _T_786 = _T_401 ? 1'h0 : _T_785; // @[Lookup.scala 33:37]
  assign _T_787 = _T_399 ? 1'h0 : _T_786; // @[Lookup.scala 33:37]
  assign _T_788 = _T_397 ? 1'h0 : _T_787; // @[Lookup.scala 33:37]
  assign _T_789 = _T_395 ? 1'h0 : _T_788; // @[Lookup.scala 33:37]
  assign _T_790 = _T_393 ? 1'h0 : _T_789; // @[Lookup.scala 33:37]
  assign _T_791 = _T_391 ? 1'h0 : _T_790; // @[Lookup.scala 33:37]
  assign _T_792 = _T_389 ? 1'h0 : _T_791; // @[Lookup.scala 33:37]
  assign _T_793 = _T_387 ? 1'h0 : _T_792; // @[Lookup.scala 33:37]
  assign _T_794 = _T_385 ? 1'h0 : _T_793; // @[Lookup.scala 33:37]
  assign _T_795 = _T_383 ? 1'h0 : _T_794; // @[Lookup.scala 33:37]
  assign _T_796 = _T_381 ? 1'h0 : _T_795; // @[Lookup.scala 33:37]
  assign _T_797 = _T_379 | _T_796; // @[Lookup.scala 33:37]
  assign _T_798 = _T_377 | _T_797; // @[Lookup.scala 33:37]
  assign _T_799 = _T_375 | _T_798; // @[Lookup.scala 33:37]
  assign _T_800 = _T_373 ? 1'h0 : _T_799; // @[Lookup.scala 33:37]
  assign _T_801 = _T_371 ? 1'h0 : _T_800; // @[Lookup.scala 33:37]
  assign _T_802 = _T_369 ? 1'h0 : _T_801; // @[Lookup.scala 33:37]
  assign _T_803 = _T_367 ? 1'h0 : _T_802; // @[Lookup.scala 33:37]
  assign _T_804 = _T_365 ? 1'h0 : _T_803; // @[Lookup.scala 33:37]
  assign _T_805 = _T_363 | _T_804; // @[Lookup.scala 33:37]
  assign _T_806 = _T_361 | _T_805; // @[Lookup.scala 33:37]
  assign _T_807 = _T_359 | _T_806; // @[Lookup.scala 33:37]
  assign _T_808 = _T_357 | _T_807; // @[Lookup.scala 33:37]
  assign _T_809 = _T_355 | _T_808; // @[Lookup.scala 33:37]
  assign _T_810 = _T_353 | _T_809; // @[Lookup.scala 33:37]
  assign _T_811 = _T_351 ? 1'h0 : _T_810; // @[Lookup.scala 33:37]
  assign _T_812 = _T_349 ? 1'h0 : _T_811; // @[Lookup.scala 33:37]
  assign _T_813 = _T_347 | _T_812; // @[Lookup.scala 33:37]
  assign _T_814 = _T_345 | _T_813; // @[Lookup.scala 33:37]
  assign _T_815 = _T_343 | _T_814; // @[Lookup.scala 33:37]
  assign _T_816 = _T_341 | _T_815; // @[Lookup.scala 33:37]
  assign _T_817 = _T_339 | _T_816; // @[Lookup.scala 33:37]
  assign _T_818 = _T_337 | _T_817; // @[Lookup.scala 33:37]
  assign _T_819 = _T_335 | _T_818; // @[Lookup.scala 33:37]
  assign _T_820 = _T_333 | _T_819; // @[Lookup.scala 33:37]
  assign _T_821 = _T_331 | _T_820; // @[Lookup.scala 33:37]
  assign _T_822 = _T_329 | _T_821; // @[Lookup.scala 33:37]
  assign _T_823 = _T_327 | _T_822; // @[Lookup.scala 33:37]
  assign _T_824 = _T_325 | _T_823; // @[Lookup.scala 33:37]
  assign _T_825 = _T_323 | _T_824; // @[Lookup.scala 33:37]
  assign _T_826 = _T_321 | _T_825; // @[Lookup.scala 33:37]
  assign _T_827 = _T_319 | _T_826; // @[Lookup.scala 33:37]
  assign _T_828 = _T_317 | _T_827; // @[Lookup.scala 33:37]
  assign _T_829 = _T_315 | _T_828; // @[Lookup.scala 33:37]
  assign _T_830 = _T_313 | _T_829; // @[Lookup.scala 33:37]
  assign _T_831 = _T_311 ? 1'h0 : _T_830; // @[Lookup.scala 33:37]
  assign _T_832 = _T_309 ? 1'h0 : _T_831; // @[Lookup.scala 33:37]
  assign _T_833 = _T_307 ? 1'h0 : _T_832; // @[Lookup.scala 33:37]
  assign _T_834 = _T_305 ? 1'h0 : _T_833; // @[Lookup.scala 33:37]
  assign _T_835 = _T_303 ? 1'h0 : _T_834; // @[Lookup.scala 33:37]
  assign _T_836 = _T_301 ? 1'h0 : _T_835; // @[Lookup.scala 33:37]
  assign _T_837 = _T_299 ? 1'h0 : _T_836; // @[Lookup.scala 33:37]
  assign _T_838 = _T_297 ? 1'h0 : _T_837; // @[Lookup.scala 33:37]
  assign _T_839 = _T_295 ? 1'h0 : _T_838; // @[Lookup.scala 33:37]
  assign _T_840 = _T_293 ? 1'h0 : _T_839; // @[Lookup.scala 33:37]
  assign _T_841 = _T_291 ? 1'h0 : _T_840; // @[Lookup.scala 33:37]
  assign _T_911 = _T_427 ? io_reg1_o : 32'h0; // @[Lookup.scala 33:37]
  assign _T_912 = _T_425 ? io_reg1_o : _T_911; // @[Lookup.scala 33:37]
  assign _T_913 = _T_423 ? io_reg1_o : _T_912; // @[Lookup.scala 33:37]
  assign _T_914 = _T_421 ? io_reg1_o : _T_913; // @[Lookup.scala 33:37]
  assign _T_915 = _T_419 ? io_reg1_o : _T_914; // @[Lookup.scala 33:37]
  assign _T_916 = _T_417 ? io_reg1_o : _T_915; // @[Lookup.scala 33:37]
  assign _T_917 = _T_415 ? io_reg1_o : _T_916; // @[Lookup.scala 33:37]
  assign _T_918 = _T_413 ? io_reg1_o : _T_917; // @[Lookup.scala 33:37]
  assign _T_919 = _T_411 ? io_reg1_o : _T_918; // @[Lookup.scala 33:37]
  assign _T_920 = _T_409 ? io_reg1_o : _T_919; // @[Lookup.scala 33:37]
  assign _T_921 = _T_407 ? io_reg1_o : _T_920; // @[Lookup.scala 33:37]
  assign _T_922 = _T_405 ? 32'h0 : _T_921; // @[Lookup.scala 33:37]
  assign _T_923 = _T_403 ? 32'h0 : _T_922; // @[Lookup.scala 33:37]
  assign _T_924 = _T_401 ? 32'h0 : _T_923; // @[Lookup.scala 33:37]
  assign _T_925 = _T_399 ? 32'h0 : _T_924; // @[Lookup.scala 33:37]
  assign _T_926 = _T_397 ? 32'h0 : _T_925; // @[Lookup.scala 33:37]
  assign _T_927 = _T_395 ? 32'h0 : _T_926; // @[Lookup.scala 33:37]
  assign _T_928 = _T_393 ? 32'h0 : _T_927; // @[Lookup.scala 33:37]
  assign _T_929 = _T_391 ? 32'h0 : _T_928; // @[Lookup.scala 33:37]
  assign _T_930 = _T_389 ? 32'h0 : _T_929; // @[Lookup.scala 33:37]
  assign _T_931 = _T_387 ? 32'h0 : _T_930; // @[Lookup.scala 33:37]
  assign _T_932 = _T_385 ? 32'h0 : _T_931; // @[Lookup.scala 33:37]
  assign _T_933 = _T_383 ? 32'h0 : _T_932; // @[Lookup.scala 33:37]
  assign _T_934 = _T_381 ? 32'h0 : _T_933; // @[Lookup.scala 33:37]
  assign _T_935 = _T_379 ? _T_250 : _T_934; // @[Lookup.scala 33:37]
  assign _T_936 = _T_377 ? _T_250 : _T_935; // @[Lookup.scala 33:37]
  assign _T_937 = _T_375 ? _T_250 : _T_936; // @[Lookup.scala 33:37]
  assign _T_938 = _T_373 ? _T_240 : _T_937; // @[Lookup.scala 33:37]
  assign _T_939 = _T_371 ? _T_240 : _T_938; // @[Lookup.scala 33:37]
  assign _T_940 = _T_369 ? _T_240 : _T_939; // @[Lookup.scala 33:37]
  assign _T_941 = _T_367 ? _T_240 : _T_940; // @[Lookup.scala 33:37]
  assign _T_942 = _T_365 ? _T_240 : _T_941; // @[Lookup.scala 33:37]
  assign _T_943 = _T_363 ? 32'h0 : _T_942; // @[Lookup.scala 33:37]
  assign _T_944 = _T_361 ? 32'h0 : _T_943; // @[Lookup.scala 33:37]
  assign _T_945 = _T_359 ? 32'h0 : _T_944; // @[Lookup.scala 33:37]
  assign _T_946 = _T_357 ? 32'h0 : _T_945; // @[Lookup.scala 33:37]
  assign _T_947 = _T_355 ? 32'h0 : _T_946; // @[Lookup.scala 33:37]
  assign _T_948 = _T_353 ? 32'h0 : _T_947; // @[Lookup.scala 33:37]
  assign _T_949 = _T_351 ? 32'h0 : _T_948; // @[Lookup.scala 33:37]
  assign _T_950 = _T_349 ? 32'h0 : _T_949; // @[Lookup.scala 33:37]
  assign _T_951 = _T_347 ? 32'h0 : _T_950; // @[Lookup.scala 33:37]
  assign _T_952 = _T_345 ? 32'h0 : _T_951; // @[Lookup.scala 33:37]
  assign _T_953 = _T_343 ? 32'h0 : _T_952; // @[Lookup.scala 33:37]
  assign _T_954 = _T_341 ? 32'h0 : _T_953; // @[Lookup.scala 33:37]
  assign _T_955 = _T_339 ? 32'h0 : _T_954; // @[Lookup.scala 33:37]
  assign _T_956 = _T_337 ? 32'h0 : _T_955; // @[Lookup.scala 33:37]
  assign _T_957 = _T_335 ? 32'h0 : _T_956; // @[Lookup.scala 33:37]
  assign _T_958 = _T_333 ? 32'h0 : _T_957; // @[Lookup.scala 33:37]
  assign _T_959 = _T_331 ? 32'h0 : _T_958; // @[Lookup.scala 33:37]
  assign _T_960 = _T_329 ? 32'h0 : _T_959; // @[Lookup.scala 33:37]
  assign _T_961 = _T_327 ? 32'h0 : _T_960; // @[Lookup.scala 33:37]
  assign _T_962 = _T_325 ? 32'h0 : _T_961; // @[Lookup.scala 33:37]
  assign _T_963 = _T_323 ? 32'h0 : _T_962; // @[Lookup.scala 33:37]
  assign _T_964 = _T_321 ? 32'h0 : _T_963; // @[Lookup.scala 33:37]
  assign _T_965 = _T_319 ? 32'h0 : _T_964; // @[Lookup.scala 33:37]
  assign _T_966 = _T_317 ? 32'h0 : _T_965; // @[Lookup.scala 33:37]
  assign _T_967 = _T_315 ? 32'h0 : _T_966; // @[Lookup.scala 33:37]
  assign _T_968 = _T_313 ? 32'h0 : _T_967; // @[Lookup.scala 33:37]
  assign _T_969 = _T_311 ? 32'h0 : _T_968; // @[Lookup.scala 33:37]
  assign _T_970 = _T_309 ? 32'h0 : _T_969; // @[Lookup.scala 33:37]
  assign _T_971 = _T_307 ? 32'h0 : _T_970; // @[Lookup.scala 33:37]
  assign _T_972 = _T_305 ? 32'h0 : _T_971; // @[Lookup.scala 33:37]
  assign _T_973 = _T_303 ? 32'h0 : _T_972; // @[Lookup.scala 33:37]
  assign _T_974 = _T_301 ? 32'h0 : _T_973; // @[Lookup.scala 33:37]
  assign _T_975 = _T_299 ? 32'h0 : _T_974; // @[Lookup.scala 33:37]
  assign _T_976 = _T_297 ? 32'h0 : _T_975; // @[Lookup.scala 33:37]
  assign _T_977 = _T_295 ? 32'h0 : _T_976; // @[Lookup.scala 33:37]
  assign _T_978 = _T_293 ? 32'h0 : _T_977; // @[Lookup.scala 33:37]
  assign _T_979 = _T_291 ? 32'h0 : _T_978; // @[Lookup.scala 33:37]
  assign _T_1012 = _T_363 ? _T_234 : 32'h0; // @[Lookup.scala 33:37]
  assign _T_1013 = _T_361 ? _T_222 : _T_1012; // @[Lookup.scala 33:37]
  assign _T_1014 = _T_359 ? _T_212 : _T_1013; // @[Lookup.scala 33:37]
  assign _T_1015 = _T_357 ? _T_200 : _T_1014; // @[Lookup.scala 33:37]
  assign _T_1016 = _T_355 ? _T_190 : _T_1015; // @[Lookup.scala 33:37]
  assign _T_1017 = _T_353 ? _T_182 : _T_1016; // @[Lookup.scala 33:37]
  assign _T_1018 = _T_351 ? _T_178 : _T_1017; // @[Lookup.scala 33:37]
  assign _T_1019 = _T_349 ? _T_174 : _T_1018; // @[Lookup.scala 33:37]
  assign _T_1020 = _T_347 ? 32'h0 : _T_1019; // @[Lookup.scala 33:37]
  assign _T_1021 = _T_345 ? 32'h0 : _T_1020; // @[Lookup.scala 33:37]
  assign _T_1022 = _T_343 ? 32'h0 : _T_1021; // @[Lookup.scala 33:37]
  assign _T_1023 = _T_341 ? 32'h0 : _T_1022; // @[Lookup.scala 33:37]
  assign _T_1024 = _T_339 ? 32'h0 : _T_1023; // @[Lookup.scala 33:37]
  assign _T_1025 = _T_337 ? 32'h0 : _T_1024; // @[Lookup.scala 33:37]
  assign _T_1026 = _T_335 ? 32'h0 : _T_1025; // @[Lookup.scala 33:37]
  assign _T_1027 = _T_333 ? 32'h0 : _T_1026; // @[Lookup.scala 33:37]
  assign _T_1028 = _T_331 ? 32'h0 : _T_1027; // @[Lookup.scala 33:37]
  assign _T_1029 = _T_329 ? 32'h0 : _T_1028; // @[Lookup.scala 33:37]
  assign _T_1030 = _T_327 ? 32'h0 : _T_1029; // @[Lookup.scala 33:37]
  assign _T_1031 = _T_325 ? 32'h0 : _T_1030; // @[Lookup.scala 33:37]
  assign _T_1032 = _T_323 ? 32'h0 : _T_1031; // @[Lookup.scala 33:37]
  assign _T_1033 = _T_321 ? 32'h0 : _T_1032; // @[Lookup.scala 33:37]
  assign _T_1034 = _T_319 ? 32'h0 : _T_1033; // @[Lookup.scala 33:37]
  assign _T_1035 = _T_317 ? 32'h0 : _T_1034; // @[Lookup.scala 33:37]
  assign _T_1036 = _T_315 ? 32'h0 : _T_1035; // @[Lookup.scala 33:37]
  assign _T_1037 = _T_313 ? 32'h0 : _T_1036; // @[Lookup.scala 33:37]
  assign _T_1038 = _T_311 ? 32'h0 : _T_1037; // @[Lookup.scala 33:37]
  assign _T_1039 = _T_309 ? 32'h0 : _T_1038; // @[Lookup.scala 33:37]
  assign _T_1040 = _T_307 ? 32'h0 : _T_1039; // @[Lookup.scala 33:37]
  assign _T_1041 = _T_305 ? 32'h0 : _T_1040; // @[Lookup.scala 33:37]
  assign _T_1042 = _T_303 ? 32'h0 : _T_1041; // @[Lookup.scala 33:37]
  assign _T_1043 = _T_301 ? 32'h0 : _T_1042; // @[Lookup.scala 33:37]
  assign _T_1044 = _T_299 ? 32'h0 : _T_1043; // @[Lookup.scala 33:37]
  assign _T_1045 = _T_297 ? 32'h0 : _T_1044; // @[Lookup.scala 33:37]
  assign _T_1046 = _T_295 ? 32'h0 : _T_1045; // @[Lookup.scala 33:37]
  assign _T_1047 = _T_293 ? 32'h0 : _T_1046; // @[Lookup.scala 33:37]
  assign _T_1048 = _T_291 ? 32'h0 : _T_1047; // @[Lookup.scala 33:37]
  assign _T_1081 = _T_363 & _T_231; // @[Lookup.scala 33:37]
  assign _T_1082 = _T_361 ? _T_219 : _T_1081; // @[Lookup.scala 33:37]
  assign _T_1083 = _T_359 ? _T_209 : _T_1082; // @[Lookup.scala 33:37]
  assign _T_1084 = _T_357 ? _T_197 : _T_1083; // @[Lookup.scala 33:37]
  assign _T_1085 = _T_355 ? _T_187 : _T_1084; // @[Lookup.scala 33:37]
  assign _T_1086 = _T_353 ? _T_179 : _T_1085; // @[Lookup.scala 33:37]
  assign _T_1087 = _T_351 | _T_1086; // @[Lookup.scala 33:37]
  assign _T_1088 = _T_349 | _T_1087; // @[Lookup.scala 33:37]
  assign _T_1089 = _T_347 ? 1'h0 : _T_1088; // @[Lookup.scala 33:37]
  assign _T_1090 = _T_345 ? 1'h0 : _T_1089; // @[Lookup.scala 33:37]
  assign _T_1091 = _T_343 ? 1'h0 : _T_1090; // @[Lookup.scala 33:37]
  assign _T_1092 = _T_341 ? 1'h0 : _T_1091; // @[Lookup.scala 33:37]
  assign _T_1093 = _T_339 ? 1'h0 : _T_1092; // @[Lookup.scala 33:37]
  assign _T_1094 = _T_337 ? 1'h0 : _T_1093; // @[Lookup.scala 33:37]
  assign _T_1095 = _T_335 ? 1'h0 : _T_1094; // @[Lookup.scala 33:37]
  assign _T_1096 = _T_333 ? 1'h0 : _T_1095; // @[Lookup.scala 33:37]
  assign _T_1097 = _T_331 ? 1'h0 : _T_1096; // @[Lookup.scala 33:37]
  assign _T_1098 = _T_329 ? 1'h0 : _T_1097; // @[Lookup.scala 33:37]
  assign _T_1099 = _T_327 ? 1'h0 : _T_1098; // @[Lookup.scala 33:37]
  assign _T_1100 = _T_325 ? 1'h0 : _T_1099; // @[Lookup.scala 33:37]
  assign _T_1101 = _T_323 ? 1'h0 : _T_1100; // @[Lookup.scala 33:37]
  assign _T_1102 = _T_321 ? 1'h0 : _T_1101; // @[Lookup.scala 33:37]
  assign _T_1103 = _T_319 ? 1'h0 : _T_1102; // @[Lookup.scala 33:37]
  assign _T_1104 = _T_317 ? 1'h0 : _T_1103; // @[Lookup.scala 33:37]
  assign _T_1105 = _T_315 ? 1'h0 : _T_1104; // @[Lookup.scala 33:37]
  assign _T_1106 = _T_313 ? 1'h0 : _T_1105; // @[Lookup.scala 33:37]
  assign _T_1107 = _T_311 ? 1'h0 : _T_1106; // @[Lookup.scala 33:37]
  assign _T_1108 = _T_309 ? 1'h0 : _T_1107; // @[Lookup.scala 33:37]
  assign _T_1109 = _T_307 ? 1'h0 : _T_1108; // @[Lookup.scala 33:37]
  assign _T_1110 = _T_305 ? 1'h0 : _T_1109; // @[Lookup.scala 33:37]
  assign _T_1111 = _T_303 ? 1'h0 : _T_1110; // @[Lookup.scala 33:37]
  assign _T_1112 = _T_301 ? 1'h0 : _T_1111; // @[Lookup.scala 33:37]
  assign _T_1113 = _T_299 ? 1'h0 : _T_1112; // @[Lookup.scala 33:37]
  assign _T_1114 = _T_297 ? 1'h0 : _T_1113; // @[Lookup.scala 33:37]
  assign _T_1115 = _T_295 ? 1'h0 : _T_1114; // @[Lookup.scala 33:37]
  assign _T_1116 = _T_293 ? 1'h0 : _T_1115; // @[Lookup.scala 33:37]
  assign _T_1117 = _T_291 ? 1'h0 : _T_1116; // @[Lookup.scala 33:37]
  assign _T_1481 = _T_391 & _T_274; // @[Lookup.scala 33:37]
  assign _T_1554 = _T_383 & _T_266; // @[Lookup.scala 33:37]
  assign _T_1613 = _T_403 | _T_405; // @[Lookup.scala 33:37]
  assign _T_1614 = _T_401 ? _T_278 : _T_1613; // @[Lookup.scala 33:37]
  assign _T_1615 = _T_399 | _T_1614; // @[Lookup.scala 33:37]
  assign _T_1616 = _T_397 | _T_1615; // @[Lookup.scala 33:37]
  assign _T_1617 = _T_395 ? _T_278 : _T_1616; // @[Lookup.scala 33:37]
  assign _T_1618 = _T_393 ? 1'h0 : _T_1617; // @[Lookup.scala 33:37]
  assign _T_1619 = _T_391 ? 1'h0 : _T_1618; // @[Lookup.scala 33:37]
  assign _T_1620 = _T_389 ? 1'h0 : _T_1619; // @[Lookup.scala 33:37]
  assign _T_1621 = _T_387 ? 1'h0 : _T_1620; // @[Lookup.scala 33:37]
  assign _T_1622 = _T_385 ? 1'h0 : _T_1621; // @[Lookup.scala 33:37]
  assign _T_1623 = _T_383 ? 1'h0 : _T_1622; // @[Lookup.scala 33:37]
  assign _T_1624 = _T_381 ? 1'h0 : _T_1623; // @[Lookup.scala 33:37]
  assign _T_1625 = _T_379 ? 1'h0 : _T_1624; // @[Lookup.scala 33:37]
  assign _T_1626 = _T_377 ? 1'h0 : _T_1625; // @[Lookup.scala 33:37]
  assign _T_1627 = _T_375 ? 1'h0 : _T_1626; // @[Lookup.scala 33:37]
  assign _T_1628 = _T_373 ? 1'h0 : _T_1627; // @[Lookup.scala 33:37]
  assign _T_1629 = _T_371 ? 1'h0 : _T_1628; // @[Lookup.scala 33:37]
  assign _T_1630 = _T_369 ? 1'h0 : _T_1629; // @[Lookup.scala 33:37]
  assign _T_1631 = _T_367 ? 1'h0 : _T_1630; // @[Lookup.scala 33:37]
  assign _T_1632 = _T_365 ? 1'h0 : _T_1631; // @[Lookup.scala 33:37]
  assign _T_1633 = _T_363 ? 1'h0 : _T_1632; // @[Lookup.scala 33:37]
  assign _T_1634 = _T_361 ? 1'h0 : _T_1633; // @[Lookup.scala 33:37]
  assign _T_1635 = _T_359 ? 1'h0 : _T_1634; // @[Lookup.scala 33:37]
  assign _T_1636 = _T_357 ? 1'h0 : _T_1635; // @[Lookup.scala 33:37]
  assign _T_1637 = _T_355 ? 1'h0 : _T_1636; // @[Lookup.scala 33:37]
  assign _T_1638 = _T_353 ? 1'h0 : _T_1637; // @[Lookup.scala 33:37]
  assign _T_1639 = _T_351 ? 1'h0 : _T_1638; // @[Lookup.scala 33:37]
  assign _T_1640 = _T_349 ? 1'h0 : _T_1639; // @[Lookup.scala 33:37]
  assign _T_1641 = _T_347 ? 1'h0 : _T_1640; // @[Lookup.scala 33:37]
  assign _T_1642 = _T_345 ? 1'h0 : _T_1641; // @[Lookup.scala 33:37]
  assign _T_1643 = _T_343 ? 1'h0 : _T_1642; // @[Lookup.scala 33:37]
  assign _T_1644 = _T_341 ? 1'h0 : _T_1643; // @[Lookup.scala 33:37]
  assign _T_1645 = _T_339 ? 1'h0 : _T_1644; // @[Lookup.scala 33:37]
  assign _T_1646 = _T_337 ? 1'h0 : _T_1645; // @[Lookup.scala 33:37]
  assign _T_1647 = _T_335 ? 1'h0 : _T_1646; // @[Lookup.scala 33:37]
  assign _T_1648 = _T_333 ? 1'h0 : _T_1647; // @[Lookup.scala 33:37]
  assign _T_1649 = _T_331 ? 1'h0 : _T_1648; // @[Lookup.scala 33:37]
  assign _T_1650 = _T_329 ? 1'h0 : _T_1649; // @[Lookup.scala 33:37]
  assign _T_1651 = _T_327 ? 1'h0 : _T_1650; // @[Lookup.scala 33:37]
  assign _T_1652 = _T_325 ? 1'h0 : _T_1651; // @[Lookup.scala 33:37]
  assign _T_1653 = _T_323 ? 1'h0 : _T_1652; // @[Lookup.scala 33:37]
  assign _T_1654 = _T_321 ? 1'h0 : _T_1653; // @[Lookup.scala 33:37]
  assign _T_1655 = _T_319 ? 1'h0 : _T_1654; // @[Lookup.scala 33:37]
  assign _T_1656 = _T_317 ? 1'h0 : _T_1655; // @[Lookup.scala 33:37]
  assign _T_1657 = _T_315 ? 1'h0 : _T_1656; // @[Lookup.scala 33:37]
  assign _T_1658 = _T_313 ? 1'h0 : _T_1657; // @[Lookup.scala 33:37]
  assign _T_1659 = _T_311 ? 1'h0 : _T_1658; // @[Lookup.scala 33:37]
  assign _T_1660 = _T_309 ? 1'h0 : _T_1659; // @[Lookup.scala 33:37]
  assign _T_1661 = _T_307 ? 1'h0 : _T_1660; // @[Lookup.scala 33:37]
  assign _T_1662 = _T_305 ? 1'h0 : _T_1661; // @[Lookup.scala 33:37]
  assign _T_1663 = _T_303 ? 1'h0 : _T_1662; // @[Lookup.scala 33:37]
  assign _T_1664 = _T_301 ? 1'h0 : _T_1663; // @[Lookup.scala 33:37]
  assign _T_1665 = _T_299 ? 1'h0 : _T_1664; // @[Lookup.scala 33:37]
  assign _T_1666 = _T_297 ? 1'h0 : _T_1665; // @[Lookup.scala 33:37]
  assign _T_1667 = _T_295 ? 1'h0 : _T_1666; // @[Lookup.scala 33:37]
  assign _T_1668 = _T_293 ? 1'h0 : _T_1667; // @[Lookup.scala 33:37]
  assign _T_1669 = _T_291 ? 1'h0 : _T_1668; // @[Lookup.scala 33:37]
  assign _T_1681 = _T_405 & _T_280; // @[Lookup.scala 33:37]
  assign _T_1682 = _T_403 ? _T_280 : _T_1681; // @[Lookup.scala 33:37]
  assign _T_1683 = _T_401 | _T_1682; // @[Lookup.scala 33:37]
  assign _T_1684 = _T_399 ? _T_280 : _T_1683; // @[Lookup.scala 33:37]
  assign _T_1685 = _T_397 ? _T_280 : _T_1684; // @[Lookup.scala 33:37]
  assign _T_1686 = _T_395 | _T_1685; // @[Lookup.scala 33:37]
  assign _T_1687 = _T_393 ? 1'h0 : _T_1686; // @[Lookup.scala 33:37]
  assign _T_1688 = _T_391 ? 1'h0 : _T_1687; // @[Lookup.scala 33:37]
  assign _T_1689 = _T_389 ? 1'h0 : _T_1688; // @[Lookup.scala 33:37]
  assign _T_1690 = _T_387 ? 1'h0 : _T_1689; // @[Lookup.scala 33:37]
  assign _T_1691 = _T_385 ? 1'h0 : _T_1690; // @[Lookup.scala 33:37]
  assign _T_1692 = _T_383 ? 1'h0 : _T_1691; // @[Lookup.scala 33:37]
  assign _T_1693 = _T_381 ? 1'h0 : _T_1692; // @[Lookup.scala 33:37]
  assign _T_1694 = _T_379 ? 1'h0 : _T_1693; // @[Lookup.scala 33:37]
  assign _T_1695 = _T_377 ? 1'h0 : _T_1694; // @[Lookup.scala 33:37]
  assign _T_1696 = _T_375 ? 1'h0 : _T_1695; // @[Lookup.scala 33:37]
  assign _T_1697 = _T_373 ? 1'h0 : _T_1696; // @[Lookup.scala 33:37]
  assign _T_1698 = _T_371 ? 1'h0 : _T_1697; // @[Lookup.scala 33:37]
  assign _T_1699 = _T_369 ? 1'h0 : _T_1698; // @[Lookup.scala 33:37]
  assign _T_1700 = _T_367 ? 1'h0 : _T_1699; // @[Lookup.scala 33:37]
  assign _T_1701 = _T_365 ? 1'h0 : _T_1700; // @[Lookup.scala 33:37]
  assign _T_1702 = _T_363 ? 1'h0 : _T_1701; // @[Lookup.scala 33:37]
  assign _T_1703 = _T_361 ? 1'h0 : _T_1702; // @[Lookup.scala 33:37]
  assign _T_1704 = _T_359 ? 1'h0 : _T_1703; // @[Lookup.scala 33:37]
  assign _T_1705 = _T_357 ? 1'h0 : _T_1704; // @[Lookup.scala 33:37]
  assign _T_1706 = _T_355 ? 1'h0 : _T_1705; // @[Lookup.scala 33:37]
  assign _T_1707 = _T_353 ? 1'h0 : _T_1706; // @[Lookup.scala 33:37]
  assign _T_1708 = _T_351 ? 1'h0 : _T_1707; // @[Lookup.scala 33:37]
  assign _T_1709 = _T_349 ? 1'h0 : _T_1708; // @[Lookup.scala 33:37]
  assign _T_1710 = _T_347 ? 1'h0 : _T_1709; // @[Lookup.scala 33:37]
  assign _T_1711 = _T_345 ? 1'h0 : _T_1710; // @[Lookup.scala 33:37]
  assign _T_1712 = _T_343 ? 1'h0 : _T_1711; // @[Lookup.scala 33:37]
  assign _T_1713 = _T_341 ? 1'h0 : _T_1712; // @[Lookup.scala 33:37]
  assign _T_1714 = _T_339 ? 1'h0 : _T_1713; // @[Lookup.scala 33:37]
  assign _T_1715 = _T_337 ? 1'h0 : _T_1714; // @[Lookup.scala 33:37]
  assign _T_1716 = _T_335 ? 1'h0 : _T_1715; // @[Lookup.scala 33:37]
  assign _T_1717 = _T_333 ? 1'h0 : _T_1716; // @[Lookup.scala 33:37]
  assign _T_1718 = _T_331 ? 1'h0 : _T_1717; // @[Lookup.scala 33:37]
  assign _T_1719 = _T_329 ? 1'h0 : _T_1718; // @[Lookup.scala 33:37]
  assign _T_1720 = _T_327 ? 1'h0 : _T_1719; // @[Lookup.scala 33:37]
  assign _T_1721 = _T_325 ? 1'h0 : _T_1720; // @[Lookup.scala 33:37]
  assign _T_1722 = _T_323 ? 1'h0 : _T_1721; // @[Lookup.scala 33:37]
  assign _T_1723 = _T_321 ? 1'h0 : _T_1722; // @[Lookup.scala 33:37]
  assign _T_1724 = _T_319 ? 1'h0 : _T_1723; // @[Lookup.scala 33:37]
  assign _T_1725 = _T_317 ? 1'h0 : _T_1724; // @[Lookup.scala 33:37]
  assign _T_1726 = _T_315 ? 1'h0 : _T_1725; // @[Lookup.scala 33:37]
  assign _T_1727 = _T_313 ? 1'h0 : _T_1726; // @[Lookup.scala 33:37]
  assign _T_1728 = _T_311 ? 1'h0 : _T_1727; // @[Lookup.scala 33:37]
  assign _T_1729 = _T_309 ? 1'h0 : _T_1728; // @[Lookup.scala 33:37]
  assign _T_1730 = _T_307 ? 1'h0 : _T_1729; // @[Lookup.scala 33:37]
  assign _T_1731 = _T_305 ? 1'h0 : _T_1730; // @[Lookup.scala 33:37]
  assign _T_1732 = _T_303 ? 1'h0 : _T_1731; // @[Lookup.scala 33:37]
  assign _T_1733 = _T_301 ? 1'h0 : _T_1732; // @[Lookup.scala 33:37]
  assign _T_1734 = _T_299 ? 1'h0 : _T_1733; // @[Lookup.scala 33:37]
  assign _T_1735 = _T_297 ? 1'h0 : _T_1734; // @[Lookup.scala 33:37]
  assign _T_1736 = _T_295 ? 1'h0 : _T_1735; // @[Lookup.scala 33:37]
  assign _T_1737 = _T_293 ? 1'h0 : _T_1736; // @[Lookup.scala 33:37]
  assign _T_1738 = _T_291 ? 1'h0 : _T_1737; // @[Lookup.scala 33:37]
  assign _T_1742 = io_reg1_read_o & _T_255; // @[IDecode.scala 1016:40]
  assign _T_1745 = io_reg1_read_o & pre_inst_is_load; // @[IDecode.scala 1018:40]
  assign _T_1747 = _T_1745 & io_ex_wreg_i; // @[IDecode.scala 1018:71]
  assign _T_1748 = io_ex_wd_i == io_reg1_addr_o; // @[IDecode.scala 1018:112]
  assign _T_1749 = _T_1747 & _T_1748; // @[IDecode.scala 1018:98]
  assign _T_1752 = io_reg1_read_o & io_ex_wreg_i; // @[IDecode.scala 1021:40]
  assign _T_1754 = _T_1752 & _T_1748; // @[IDecode.scala 1021:67]
  assign _T_1757 = io_reg1_read_o & io_mem_wreg_i; // @[IDecode.scala 1023:40]
  assign _T_1758 = io_mem_wd_i == io_reg1_addr_o; // @[IDecode.scala 1023:83]
  assign _T_1759 = _T_1757 & _T_1758; // @[IDecode.scala 1023:68]
  assign _GEN_93 = io_reg1_read_o ? 32'h0 : imm; // @[IDecode.scala 1027:41]
  assign _GEN_94 = io_reg1_read_o ? io_reg1_data_i : _GEN_93; // @[IDecode.scala 1025:40]
  assign _GEN_95 = _T_1759 ? io_mem_wdata_i : _GEN_94; // @[IDecode.scala 1023:102]
  assign _GEN_96 = _T_1754 ? io_ex_wdata_i : _GEN_95; // @[IDecode.scala 1021:100]
  assign _GEN_98 = _T_1749 ? 32'h0 : _GEN_96; // @[IDecode.scala 1018:131]
  assign _GEN_99 = _T_1742 ? 32'h0 : _GEN_98; // @[IDecode.scala 1016:76]
  assign _T_1764 = io_reg2_addr_o == 5'h0; // @[IDecode.scala 1037:58]
  assign _T_1765 = io_reg2_read_o & _T_1764; // @[IDecode.scala 1037:40]
  assign _T_1768 = io_reg2_read_o & pre_inst_is_load; // @[IDecode.scala 1039:40]
  assign _T_1770 = _T_1768 & io_ex_wreg_i; // @[IDecode.scala 1039:71]
  assign _T_1771 = io_ex_wd_i == io_reg2_addr_o; // @[IDecode.scala 1039:112]
  assign _T_1772 = _T_1770 & _T_1771; // @[IDecode.scala 1039:98]
  assign _T_1775 = io_reg2_read_o & io_ex_wreg_i; // @[IDecode.scala 1042:40]
  assign _T_1777 = _T_1775 & _T_1771; // @[IDecode.scala 1042:67]
  assign _T_1780 = io_reg2_read_o & io_mem_wreg_i; // @[IDecode.scala 1044:40]
  assign _T_1781 = io_mem_wd_i == io_reg2_addr_o; // @[IDecode.scala 1044:83]
  assign _T_1782 = _T_1780 & _T_1781; // @[IDecode.scala 1044:68]
  assign _GEN_103 = io_reg2_read_o ? 32'h0 : imm; // @[IDecode.scala 1048:41]
  assign _GEN_104 = io_reg2_read_o ? io_reg2_data_i : _GEN_103; // @[IDecode.scala 1046:40]
  assign _GEN_105 = _T_1782 ? io_mem_wdata_i : _GEN_104; // @[IDecode.scala 1044:102]
  assign _GEN_106 = _T_1777 ? io_ex_wdata_i : _GEN_105; // @[IDecode.scala 1042:100]
  assign _GEN_108 = _T_1772 ? 32'h0 : _GEN_106; // @[IDecode.scala 1039:131]
  assign _GEN_109 = _T_1765 ? 32'h0 : _GEN_108; // @[IDecode.scala 1037:76]
  assign io_csr_reg_data_o = io_csr_reg_data_i; // @[IDecode.scala 198:20]
  assign io_csr_reg_read_o = _T_170 ? 1'h0 : _T_1669; // @[IDecode.scala 309:21 IDecode.scala 337:21 IDecode.scala 1008:22]
  assign io_csr_reg_we_o = _T_170 ? 1'h0 : _T_1738; // @[IDecode.scala 310:19 IDecode.scala 338:19 IDecode.scala 1009:22]
  assign io_csr_reg_addr_o = io_inst_i[31:20]; // @[IDecode.scala 194:20]
  assign io_reg1_read_o = _T_170 ? 1'h0 : _T_772; // @[IDecode.scala 291:18 IDecode.scala 319:18 IDecode.scala 990:19]
  assign io_reg2_read_o = _T_170 ? 1'h0 : _T_841; // @[IDecode.scala 292:18 IDecode.scala 320:18 IDecode.scala 991:19]
  assign io_reg1_addr_o = io_inst_i[19:15]; // @[IDecode.scala 192:17]
  assign io_reg2_addr_o = io_inst_i[24:20]; // @[IDecode.scala 193:17]
  assign io_aluop_o = _T_170 ? 8'h0 : _T_496; // @[IDecode.scala 286:14 IDecode.scala 314:14 IDecode.scala 984:19]
  assign io_alusel_o = _T_170 ? 3'h0 : _T_565; // @[IDecode.scala 287:15 IDecode.scala 315:15 IDecode.scala 985:19]
  assign io_reg1_o = io_rst_n ? _GEN_99 : 32'h0; // @[IDecode.scala 1015:15 IDecode.scala 1017:15 IDecode.scala 1020:15 IDecode.scala 1022:15 IDecode.scala 1024:15 IDecode.scala 1026:15 IDecode.scala 1028:15 IDecode.scala 1030:15]
  assign io_reg2_o = io_rst_n ? _GEN_109 : 32'h0; // @[IDecode.scala 1036:15 IDecode.scala 1038:15 IDecode.scala 1041:15 IDecode.scala 1043:15 IDecode.scala 1045:15 IDecode.scala 1047:15 IDecode.scala 1049:15 IDecode.scala 1051:15]
  assign io_mem_addr_o = _T_170 ? 32'h0 : _T_979; // @[IDecode.scala 296:17 IDecode.scala 324:17 IDecode.scala 995:19]
  assign io_wd_o = io_inst_i[11:7]; // @[IDecode.scala 196:10]
  assign io_wreg_o = _T_170 ? 1'h0 : _T_703; // @[IDecode.scala 290:13 IDecode.scala 318:13 IDecode.scala 988:19]
  assign io_inst_o = io_inst_i; // @[IDecode.scala 200:12]
  assign io_next_inst_in_delayslot_o = _T_170 ? 1'h0 : _T_1117; // @[IDecode.scala 300:31 IDecode.scala 328:31 IDecode.scala 999:32]
  assign io_branch_flag_o = _T_170 ? 1'h0 : _T_1117; // @[IDecode.scala 299:20 IDecode.scala 327:20 IDecode.scala 998:32]
  assign io_branch_target_address_o = _T_170 ? 32'h0 : _T_1048; // @[IDecode.scala 298:30 IDecode.scala 326:30 IDecode.scala 997:32]
  assign io_link_addr_o = io_pc_i + 32'h4; // @[IDecode.scala 199:17]
  assign io_is_in_delayslot_o = io_rst_n ? io_is_in_delayslot_i : 1'h0; // @[IDecode.scala 1056:26 IDecode.scala 1058:26]
  assign io_excepttype_o = io_rst_n ? _GEN_39 : 32'h0; // @[IDecode.scala 255:19 IDecode.scala 278:19]
  assign io_current_inst_address_o = io_pc_i; // @[IDecode.scala 201:28]
  assign io_not_stall_o = io_rst_n ? _GEN_6 : 1'h0; // @[IDecode.scala 258:18 IDecode.scala 261:18 IDecode.scala 279:18]
  assign io_step_o = 1'h0; // @[IDecode.scala 301:13 IDecode.scala 329:13 IDecode.scala 1000:32]
  assign io_stallreq = _T_62 | stallreq_for_csr_read_relate; // @[IDecode.scala 241:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  imm = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  imm_i_type = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  imm_s_type = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  imm_u_type = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  imm_sb_type = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  imm_uj_type = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  zimm = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  instvalid = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  stallreq_for_reg1_loadrelate = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  stallreq_for_reg2_loadrelate = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  stallreq_for_csr_write_relate = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  stallreq_for_csr_read_relate = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  pre_inst_is_load = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  excepttype_is_syscall = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  excepttype_is_break = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  excepttype_is_sret = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  excepttype_is_mret = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  excepttype_is_fence_i = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
always @(*) begin
    if (_T_170) begin
      imm <= 32'h0;
    end else if (_T_291) begin
      imm <= imm_i_type;
    end else if (_T_293) begin
      imm <= imm_i_type;
    end else if (_T_295) begin
      imm <= imm_i_type;
    end else if (_T_297) begin
      imm <= imm_i_type;
    end else if (_T_299) begin
      imm <= imm_i_type;
    end else if (_T_301) begin
      imm <= imm_i_type;
    end else if (_T_303) begin
      imm <= imm_i_type;
    end else if (_T_305) begin
      imm <= imm_i_type;
    end else if (_T_307) begin
      imm <= imm_i_type;
    end else if (_T_309) begin
      imm <= imm_u_type;
    end else if (_T_311) begin
      imm <= _T_172;
    end else if (_T_313) begin
      imm <= 32'h0;
    end else if (_T_315) begin
      imm <= 32'h0;
    end else if (_T_317) begin
      imm <= 32'h0;
    end else if (_T_319) begin
      imm <= 32'h0;
    end else if (_T_321) begin
      imm <= 32'h0;
    end else if (_T_323) begin
      imm <= 32'h0;
    end else if (_T_325) begin
      imm <= 32'h0;
    end else if (_T_327) begin
      imm <= 32'h0;
    end else if (_T_329) begin
      imm <= 32'h0;
    end else if (_T_331) begin
      imm <= 32'h0;
    end else if (_T_333) begin
      imm <= 32'h0;
    end else if (_T_335) begin
      imm <= 32'h0;
    end else if (_T_337) begin
      imm <= 32'h0;
    end else if (_T_339) begin
      imm <= 32'h0;
    end else if (_T_341) begin
      imm <= 32'h0;
    end else if (_T_343) begin
      imm <= 32'h0;
    end else if (_T_345) begin
      imm <= 32'h0;
    end else if (_T_347) begin
      imm <= 32'h0;
    end else if (_T_349) begin
      imm <= 32'h0;
    end else if (_T_351) begin
      imm <= 32'h0;
    end else if (_T_353) begin
      imm <= 32'h0;
    end else if (_T_355) begin
      imm <= 32'h0;
    end else if (_T_357) begin
      imm <= 32'h0;
    end else if (_T_359) begin
      imm <= 32'h0;
    end else if (_T_361) begin
      imm <= 32'h0;
    end else if (_T_363) begin
      imm <= 32'h0;
    end else if (_T_365) begin
      imm <= 32'h0;
    end else if (_T_367) begin
      imm <= 32'h0;
    end else if (_T_369) begin
      imm <= 32'h0;
    end else if (_T_371) begin
      imm <= 32'h0;
    end else if (_T_373) begin
      imm <= 32'h0;
    end else if (_T_375) begin
      imm <= 32'h0;
    end else if (_T_377) begin
      imm <= 32'h0;
    end else if (_T_379) begin
      imm <= 32'h0;
    end else if (_T_381) begin
      imm <= 32'h0;
    end else if (_T_383) begin
      imm <= 32'h0;
    end else if (_T_385) begin
      imm <= 32'h0;
    end else if (_T_387) begin
      imm <= 32'h0;
    end else if (_T_389) begin
      imm <= 32'h0;
    end else if (_T_391) begin
      imm <= 32'h0;
    end else if (_T_393) begin
      imm <= 32'h0;
    end else if (_T_395) begin
      imm <= 32'h0;
    end else if (_T_397) begin
      imm <= 32'h0;
    end else if (_T_399) begin
      imm <= 32'h0;
    end else if (_T_401) begin
      imm <= zimm;
    end else if (_T_403) begin
      imm <= zimm;
    end else if (_T_405) begin
      imm <= zimm;
    end else begin
      imm <= 32'h0;
    end
    imm_i_type <= {_T_12,io_inst_i[31:20]};
    imm_s_type <= {_T_19,io_inst_i[11:7]};
    imm_u_type <= {io_inst_i[31:12],12'h0};
    imm_sb_type <= {_T_35,1'h0};
    imm_uj_type <= {_T_47,1'h0};
    zimm <= {27'h0,io_inst_i[19:15]};
    if (_T_170) begin
      instvalid <= 1'h0;
    end else if (_T_291) begin
      instvalid <= 1'h0;
    end else if (_T_293) begin
      instvalid <= 1'h0;
    end else if (_T_295) begin
      instvalid <= 1'h0;
    end else if (_T_297) begin
      instvalid <= 1'h0;
    end else if (_T_299) begin
      instvalid <= 1'h0;
    end else if (_T_301) begin
      instvalid <= 1'h0;
    end else if (_T_303) begin
      instvalid <= 1'h0;
    end else if (_T_305) begin
      instvalid <= 1'h0;
    end else if (_T_307) begin
      instvalid <= 1'h0;
    end else if (_T_309) begin
      instvalid <= 1'h0;
    end else if (_T_311) begin
      instvalid <= 1'h0;
    end else if (_T_313) begin
      instvalid <= 1'h0;
    end else if (_T_315) begin
      instvalid <= 1'h0;
    end else if (_T_317) begin
      instvalid <= 1'h0;
    end else if (_T_319) begin
      instvalid <= 1'h0;
    end else if (_T_321) begin
      instvalid <= 1'h0;
    end else if (_T_323) begin
      instvalid <= 1'h0;
    end else if (_T_325) begin
      instvalid <= 1'h0;
    end else if (_T_327) begin
      instvalid <= 1'h0;
    end else if (_T_329) begin
      instvalid <= 1'h0;
    end else if (_T_331) begin
      instvalid <= 1'h0;
    end else if (_T_333) begin
      instvalid <= 1'h0;
    end else if (_T_335) begin
      instvalid <= 1'h0;
    end else if (_T_337) begin
      instvalid <= 1'h0;
    end else if (_T_339) begin
      instvalid <= 1'h0;
    end else if (_T_341) begin
      instvalid <= 1'h0;
    end else if (_T_343) begin
      instvalid <= 1'h0;
    end else if (_T_345) begin
      instvalid <= 1'h0;
    end else if (_T_347) begin
      instvalid <= 1'h0;
    end else if (_T_349) begin
      instvalid <= 1'h0;
    end else if (_T_351) begin
      instvalid <= 1'h0;
    end else if (_T_353) begin
      instvalid <= 1'h0;
    end else if (_T_355) begin
      instvalid <= 1'h0;
    end else if (_T_357) begin
      instvalid <= 1'h0;
    end else if (_T_359) begin
      instvalid <= 1'h0;
    end else if (_T_361) begin
      instvalid <= 1'h0;
    end else if (_T_363) begin
      instvalid <= 1'h0;
    end else if (_T_365) begin
      instvalid <= 1'h0;
    end else if (_T_367) begin
      instvalid <= 1'h0;
    end else if (_T_369) begin
      instvalid <= 1'h0;
    end else if (_T_371) begin
      instvalid <= 1'h0;
    end else if (_T_373) begin
      instvalid <= 1'h0;
    end else if (_T_375) begin
      instvalid <= 1'h0;
    end else if (_T_377) begin
      instvalid <= 1'h0;
    end else if (_T_379) begin
      instvalid <= 1'h0;
    end else if (_T_381) begin
      if (_T_260) begin
        instvalid <= 1'h0;
      end else begin
        instvalid <= 1'h1;
      end
    end else if (_T_383) begin
      if (_T_266) begin
        instvalid <= 1'h0;
      end else begin
        instvalid <= 1'h1;
      end
    end else if (_T_385) begin
      instvalid <= 1'h0;
    end else if (_T_387) begin
      instvalid <= 1'h0;
    end else if (_T_389) begin
      instvalid <= 1'h0;
    end else if (_T_391) begin
      if (_T_274) begin
        instvalid <= 1'h0;
      end else begin
        instvalid <= 1'h1;
      end
    end else if (_T_393) begin
      instvalid <= 1'h0;
    end else if (_T_395) begin
      instvalid <= 1'h0;
    end else if (_T_397) begin
      instvalid <= 1'h0;
    end else if (_T_399) begin
      instvalid <= 1'h0;
    end else if (_T_401) begin
      instvalid <= 1'h0;
    end else if (_T_403) begin
      instvalid <= 1'h0;
    end else if (_T_405) begin
      instvalid <= 1'h0;
    end else if (_T_407) begin
      instvalid <= 1'h0;
    end else if (_T_409) begin
      instvalid <= 1'h0;
    end else if (_T_411) begin
      instvalid <= 1'h0;
    end else if (_T_413) begin
      instvalid <= 1'h0;
    end else if (_T_415) begin
      instvalid <= 1'h0;
    end else if (_T_417) begin
      instvalid <= 1'h0;
    end else if (_T_419) begin
      instvalid <= 1'h0;
    end else if (_T_421) begin
      instvalid <= 1'h0;
    end else if (_T_423) begin
      instvalid <= 1'h0;
    end else if (_T_425) begin
      instvalid <= 1'h0;
    end else if (_T_427) begin
      instvalid <= 1'h0;
    end else begin
      instvalid <= 1'h1;
    end
    if (~io_rst_n) begin
      stallreq_for_reg1_loadrelate <= 1'h0;
    end else if (_T_1742) begin
      stallreq_for_reg1_loadrelate <= 1'h0;
    end else begin
      stallreq_for_reg1_loadrelate <= _T_1749;
    end
    if (~io_rst_n) begin
      stallreq_for_reg2_loadrelate <= 1'h0;
    end else if (_T_1765) begin
      stallreq_for_reg2_loadrelate <= 1'h0;
    end else begin
      stallreq_for_reg2_loadrelate <= _T_1772;
    end
    if (_T_56) begin
      stallreq_for_csr_write_relate <= 1'h0;
    end else begin
      stallreq_for_csr_write_relate <= 1'h1;
    end
    stallreq_for_csr_read_relate <= io_csr_reg_read_o & _T_59;
    pre_inst_is_load <= _T_92 | _T_93;
    if (_T_170) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_291) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_293) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_295) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_297) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_299) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_301) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_303) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_305) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_307) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_309) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_311) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_313) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_315) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_317) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_319) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_321) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_323) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_325) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_327) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_329) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_331) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_333) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_335) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_337) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_339) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_341) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_343) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_345) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_347) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_349) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_351) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_353) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_355) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_357) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_359) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_361) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_363) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_365) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_367) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_369) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_371) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_373) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_375) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_377) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_379) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_381) begin
      excepttype_is_syscall <= 1'h0;
    end else if (_T_383) begin
      excepttype_is_syscall <= 1'h0;
    end else begin
      excepttype_is_syscall <= _T_385;
    end
    if (_T_170) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_291) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_293) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_295) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_297) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_299) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_301) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_303) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_305) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_307) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_309) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_311) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_313) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_315) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_317) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_319) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_321) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_323) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_325) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_327) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_329) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_331) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_333) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_335) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_337) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_339) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_341) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_343) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_345) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_347) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_349) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_351) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_353) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_355) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_357) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_359) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_361) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_363) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_365) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_367) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_369) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_371) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_373) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_375) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_377) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_379) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_381) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_383) begin
      excepttype_is_break <= 1'h0;
    end else if (_T_385) begin
      excepttype_is_break <= 1'h0;
    end else begin
      excepttype_is_break <= _T_387;
    end
    if (_T_170) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_291) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_293) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_295) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_297) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_299) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_301) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_303) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_305) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_307) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_309) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_311) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_313) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_315) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_317) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_319) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_321) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_323) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_325) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_327) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_329) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_331) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_333) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_335) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_337) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_339) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_341) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_343) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_345) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_347) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_349) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_351) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_353) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_355) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_357) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_359) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_361) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_363) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_365) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_367) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_369) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_371) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_373) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_375) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_377) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_379) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_381) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_383) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_385) begin
      excepttype_is_sret <= 1'h0;
    end else if (_T_387) begin
      excepttype_is_sret <= 1'h0;
    end else begin
      excepttype_is_sret <= _T_389;
    end
    if (_T_170) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_291) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_293) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_295) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_297) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_299) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_301) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_303) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_305) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_307) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_309) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_311) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_313) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_315) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_317) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_319) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_321) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_323) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_325) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_327) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_329) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_331) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_333) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_335) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_337) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_339) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_341) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_343) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_345) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_347) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_349) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_351) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_353) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_355) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_357) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_359) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_361) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_363) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_365) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_367) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_369) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_371) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_373) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_375) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_377) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_379) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_381) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_383) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_385) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_387) begin
      excepttype_is_mret <= 1'h0;
    end else if (_T_389) begin
      excepttype_is_mret <= 1'h0;
    end else begin
      excepttype_is_mret <= _T_1481;
    end
    if (_T_170) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_291) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_293) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_295) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_297) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_299) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_301) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_303) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_305) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_307) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_309) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_311) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_313) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_315) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_317) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_319) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_321) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_323) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_325) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_327) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_329) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_331) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_333) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_335) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_337) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_339) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_341) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_343) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_345) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_347) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_349) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_351) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_353) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_355) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_357) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_359) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_361) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_363) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_365) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_367) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_369) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_371) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_373) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_375) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_377) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_379) begin
      excepttype_is_fence_i <= 1'h0;
    end else if (_T_381) begin
      excepttype_is_fence_i <= 1'h0;
    end else begin
      excepttype_is_fence_i <= _T_1554;
    end
end
endmodule
