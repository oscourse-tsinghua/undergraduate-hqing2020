module IMemory(
  input         io_rst_n,
  input  [33:0] io_mem_phy_addr_i,
  input         io_data_tlb_r_exception_i,
  input         io_data_tlb_w_exception_i,
  input  [4:0]  io_wd_i,
  input         io_wreg_i,
  input  [31:0] io_wdata_i,
  input  [7:0]  io_aluop_i,
  input  [31:0] io_mem_addr_i,
  input  [31:0] io_reg2_i,
  input  [31:0] io_mem_data_i,
  input         io_LLbit_i,
  input  [33:0] io_LLbit_addr_i,
  input         io_stallreq_from_mem_i,
  input  [1:0]  io_cnt_i,
  input  [31:0] io_original_data_i,
  input         io_csr_reg_we_i,
  input  [11:0] io_csr_reg_addr_i,
  input  [31:0] io_csr_reg_data_i,
  input  [31:0] io_excepttype_i,
  input         io_is_in_delayslot_i,
  input  [31:0] io_current_inst_address_i,
  input         io_not_stall_i,
  output [4:0]  io_wd_o,
  output        io_wreg_o,
  output [31:0] io_wdata_o,
  output        io_LLbit_we_o,
  output        io_LLbit_value_o,
  output [33:0] io_LLbit_addr_o,
  output        io_stallreq,
  output [1:0]  io_cnt_o,
  output [31:0] io_original_data_o,
  output        io_csr_reg_we_o,
  output [11:0] io_csr_reg_addr_o,
  output [31:0] io_csr_reg_data_o,
  output [31:0] io_excepttype_o,
  output        io_is_in_delayslot_o,
  output [31:0] io_current_inst_address_o,
  output [31:0] io_current_data_address_o,
  output        io_not_stall_o,
  output [31:0] io_mem_addr_o,
  output [33:0] io_mem_phy_addr_o,
  output        io_mem_we_o,
  output [3:0]  io_mem_sel_o,
  output [31:0] io_mem_data_o,
  output        io_mem_ce_o
);
  reg  stallreq_from_amo; // @[IMemory.scala 89:30]
  reg [31:0] _RAND_0;
  reg [4:0] wd_o; // @[IMemory.scala 93:21]
  reg [31:0] _RAND_1;
  reg  wreg_o; // @[IMemory.scala 94:23]
  reg [31:0] _RAND_2;
  reg [31:0] wdata_o; // @[IMemory.scala 95:24]
  reg [31:0] _RAND_3;
  reg [31:0] mem_addr_o; // @[IMemory.scala 101:27]
  reg [31:0] _RAND_4;
  reg [33:0] mem_phy_addr_o; // @[IMemory.scala 102:31]
  reg [63:0] _RAND_5;
  reg  mem_we_o; // @[IMemory.scala 103:25]
  reg [31:0] _RAND_6;
  reg [3:0] mem_sel_o; // @[IMemory.scala 104:26]
  reg [31:0] _RAND_7;
  reg [31:0] mem_data_o; // @[IMemory.scala 105:27]
  reg [31:0] _RAND_8;
  reg  mem_ce_o; // @[IMemory.scala 106:25]
  reg [31:0] _RAND_9;
  reg  LLbit_we_o; // @[IMemory.scala 108:27]
  reg [31:0] _RAND_10;
  reg [33:0] LLbit_addr_o; // @[IMemory.scala 109:29]
  reg [63:0] _RAND_11;
  reg  LLbit_value_o; // @[IMemory.scala 110:30]
  reg [31:0] _RAND_12;
  reg [1:0] cnt_o; // @[IMemory.scala 112:22]
  reg [31:0] _RAND_13;
  reg [31:0] original_data_o; // @[IMemory.scala 113:32]
  reg [31:0] _RAND_14;
  wire  _T_2; // @[IMemory.scala 198:21]
  wire  _T_4; // @[IMemory.scala 211:35]
  wire [23:0] _T_7; // @[Bitwise.scala 71:12]
  wire [31:0] _T_9; // @[Cat.scala 29:58]
  wire  _T_11; // @[IMemory.scala 215:41]
  wire [23:0] _T_14; // @[Bitwise.scala 71:12]
  wire [31:0] _T_16; // @[Cat.scala 29:58]
  wire  _T_18; // @[IMemory.scala 219:41]
  wire [23:0] _T_21; // @[Bitwise.scala 71:12]
  wire [31:0] _T_23; // @[Cat.scala 29:58]
  wire  _T_25; // @[IMemory.scala 223:41]
  wire [23:0] _T_28; // @[Bitwise.scala 71:12]
  wire [31:0] _T_30; // @[Cat.scala 29:58]
  wire  _GEN_6; // @[IMemory.scala 219:59]
  wire  _GEN_10; // @[IMemory.scala 215:59]
  wire  _GEN_14; // @[IMemory.scala 211:52]
  wire [31:0] _GEN_18; // @[IMemory.scala 199:38]
  wire [33:0] _GEN_19; // @[IMemory.scala 199:38]
  wire  _GEN_21; // @[IMemory.scala 199:38]
  wire  _T_31; // @[IMemory.scala 235:27]
  wire [31:0] _T_36; // @[Cat.scala 29:58]
  wire [31:0] _T_41; // @[Cat.scala 29:58]
  wire [31:0] _T_46; // @[Cat.scala 29:58]
  wire [31:0] _T_51; // @[Cat.scala 29:58]
  wire  _T_52; // @[IMemory.scala 272:27]
  wire [15:0] _T_57; // @[Bitwise.scala 71:12]
  wire [31:0] _T_59; // @[Cat.scala 29:58]
  wire [15:0] _T_64; // @[Bitwise.scala 71:12]
  wire [31:0] _T_66; // @[Cat.scala 29:58]
  wire  _GEN_51; // @[IMemory.scala 285:52]
  wire  _T_67; // @[IMemory.scala 301:27]
  wire [31:0] _T_72; // @[Cat.scala 29:58]
  wire [31:0] _T_77; // @[Cat.scala 29:58]
  wire  _T_78; // @[IMemory.scala 330:27]
  wire [3:0] _GEN_70; // @[IMemory.scala 343:52]
  wire  _T_81; // @[IMemory.scala 355:27]
  wire  _T_84; // @[IMemory.scala 381:27]
  wire [31:0] _T_87; // @[Cat.scala 29:58]
  wire  _GEN_101; // @[IMemory.scala 382:38]
  wire  _T_96; // @[IMemory.scala 414:27]
  wire [31:0] _T_98; // @[Cat.scala 29:58]
  wire  _T_103; // @[IMemory.scala 441:27]
  wire  _T_106; // @[IMemory.scala 464:27]
  wire  _T_108; // @[IMemory.scala 467:59]
  wire  _T_109; // @[IMemory.scala 467:40]
  wire  _GEN_124; // @[IMemory.scala 467:81]
  wire  _T_112; // @[IMemory.scala 502:27]
  wire  _T_113; // @[IMemory.scala 502:64]
  wire  _T_114; // @[IMemory.scala 502:50]
  wire  _T_115; // @[IMemory.scala 502:100]
  wire  _T_116; // @[IMemory.scala 502:86]
  wire  _T_117; // @[IMemory.scala 503:18]
  wire  _T_118; // @[IMemory.scala 502:122]
  wire  _T_119; // @[IMemory.scala 503:54]
  wire  _T_120; // @[IMemory.scala 503:40]
  wire  _T_121; // @[IMemory.scala 503:89]
  wire  _T_122; // @[IMemory.scala 503:75]
  wire  _T_123; // @[IMemory.scala 504:18]
  wire  _T_124; // @[IMemory.scala 503:111]
  wire  _T_125; // @[IMemory.scala 504:54]
  wire  _T_126; // @[IMemory.scala 504:40]
  wire  _T_127; // @[IMemory.scala 504:91]
  wire  _T_128; // @[IMemory.scala 504:77]
  wire  _T_129; // @[IMemory.scala 506:38]
  wire  _T_130; // @[IMemory.scala 508:27]
  wire  _T_135; // @[IMemory.scala 530:27]
  wire [31:0] _T_139; // @[IMemory.scala 542:92]
  wire [31:0] _T_141; // @[IMemory.scala 543:92]
  wire [31:0] _T_143; // @[IMemory.scala 544:92]
  wire [31:0] _T_145; // @[IMemory.scala 545:92]
  wire  _T_149; // @[IMemory.scala 546:103]
  wire  _T_154; // @[IMemory.scala 547:103]
  wire  _T_157; // @[IMemory.scala 548:96]
  wire  _T_160; // @[IMemory.scala 549:96]
  wire  _GEN_173; // @[IMemory.scala 508:40]
  wire  _GEN_176; // @[IMemory.scala 508:40]
  wire  _GEN_177; // @[IMemory.scala 508:40]
  wire  _GEN_180; // @[IMemory.scala 508:40]
  wire  _GEN_188; // @[IMemory.scala 506:66]
  wire  _GEN_191; // @[IMemory.scala 506:66]
  wire  _GEN_192; // @[IMemory.scala 506:66]
  wire  _GEN_195; // @[IMemory.scala 506:66]
  wire  _GEN_203; // @[IMemory.scala 504:114]
  wire  _GEN_206; // @[IMemory.scala 504:114]
  wire  _GEN_207; // @[IMemory.scala 504:114]
  wire  _GEN_210; // @[IMemory.scala 504:114]
  wire  _GEN_312; // @[IMemory.scala 355:43]
  wire [31:0] _GEN_479; // @[IMemory.scala 616:28]
  assign _T_2 = io_aluop_i == 8'he0; // @[IMemory.scala 198:21]
  assign _T_4 = io_mem_addr_i[1:0] == 2'h0; // @[IMemory.scala 211:35]
  assign _T_7 = io_mem_data_i[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 71:12]
  assign _T_9 = {_T_7,io_mem_data_i[7:0]}; // @[Cat.scala 29:58]
  assign _T_11 = io_mem_addr_i[1:0] == 2'h1; // @[IMemory.scala 215:41]
  assign _T_14 = io_mem_data_i[15] ? 24'hffffff : 24'h0; // @[Bitwise.scala 71:12]
  assign _T_16 = {_T_14,io_mem_data_i[15:8]}; // @[Cat.scala 29:58]
  assign _T_18 = io_mem_addr_i[1:0] == 2'h2; // @[IMemory.scala 219:41]
  assign _T_21 = io_mem_data_i[23] ? 24'hffffff : 24'h0; // @[Bitwise.scala 71:12]
  assign _T_23 = {_T_21,io_mem_data_i[23:16]}; // @[Cat.scala 29:58]
  assign _T_25 = io_mem_addr_i[1:0] == 2'h3; // @[IMemory.scala 223:41]
  assign _T_28 = io_mem_data_i[31] ? 24'hffffff : 24'h0; // @[Bitwise.scala 71:12]
  assign _T_30 = {_T_28,io_mem_data_i[31:24]}; // @[Cat.scala 29:58]
  assign _GEN_6 = _T_18 | _T_25; // @[IMemory.scala 219:59]
  assign _GEN_10 = _T_11 | _GEN_6; // @[IMemory.scala 215:59]
  assign _GEN_14 = _T_4 | _GEN_10; // @[IMemory.scala 211:52]
  assign _GEN_18 = io_data_tlb_r_exception_i ? 32'h0 : io_mem_addr_i; // @[IMemory.scala 199:38]
  assign _GEN_19 = io_data_tlb_r_exception_i ? 34'h0 : io_mem_phy_addr_i; // @[IMemory.scala 199:38]
  assign _GEN_21 = io_data_tlb_r_exception_i ? 1'h0 : 1'h1; // @[IMemory.scala 199:38]
  assign _T_31 = io_aluop_i == 8'he4; // @[IMemory.scala 235:27]
  assign _T_36 = {24'h0,io_mem_data_i[7:0]}; // @[Cat.scala 29:58]
  assign _T_41 = {24'h0,io_mem_data_i[15:8]}; // @[Cat.scala 29:58]
  assign _T_46 = {24'h0,io_mem_data_i[23:16]}; // @[Cat.scala 29:58]
  assign _T_51 = {24'h0,io_mem_data_i[31:24]}; // @[Cat.scala 29:58]
  assign _T_52 = io_aluop_i == 8'he1; // @[IMemory.scala 272:27]
  assign _T_57 = io_mem_data_i[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_59 = {_T_57,io_mem_data_i[15:0]}; // @[Cat.scala 29:58]
  assign _T_64 = io_mem_data_i[31] ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_66 = {_T_64,io_mem_data_i[31:16]}; // @[Cat.scala 29:58]
  assign _GEN_51 = _T_4 | _T_18; // @[IMemory.scala 285:52]
  assign _T_67 = io_aluop_i == 8'he5; // @[IMemory.scala 301:27]
  assign _T_72 = {16'h0,io_mem_data_i[15:0]}; // @[Cat.scala 29:58]
  assign _T_77 = {16'h0,io_mem_data_i[31:16]}; // @[Cat.scala 29:58]
  assign _T_78 = io_aluop_i == 8'he3; // @[IMemory.scala 330:27]
  assign _GEN_70 = _T_4 ? 4'hf : 4'h0; // @[IMemory.scala 343:52]
  assign _T_81 = io_aluop_i == 8'hf0; // @[IMemory.scala 355:27]
  assign _T_84 = io_aluop_i == 8'he8; // @[IMemory.scala 381:27]
  assign _T_87 = {io_reg2_i[7:0],io_reg2_i[7:0],io_reg2_i[7:0],io_reg2_i[7:0]}; // @[Cat.scala 29:58]
  assign _GEN_101 = io_data_tlb_w_exception_i ? 1'h0 : 1'h1; // @[IMemory.scala 382:38]
  assign _T_96 = io_aluop_i == 8'he9; // @[IMemory.scala 414:27]
  assign _T_98 = {io_reg2_i[15:0],io_reg2_i[15:0]}; // @[Cat.scala 29:58]
  assign _T_103 = io_aluop_i == 8'heb; // @[IMemory.scala 441:27]
  assign _T_106 = io_aluop_i == 8'hf8; // @[IMemory.scala 464:27]
  assign _T_108 = io_LLbit_addr_i == io_mem_phy_addr_i; // @[IMemory.scala 467:59]
  assign _T_109 = io_LLbit_i & _T_108; // @[IMemory.scala 467:40]
  assign _GEN_124 = _T_109 & _T_4; // @[IMemory.scala 467:81]
  assign _T_112 = io_aluop_i == 8'h41; // @[IMemory.scala 502:27]
  assign _T_113 = io_aluop_i == 8'h40; // @[IMemory.scala 502:64]
  assign _T_114 = _T_112 | _T_113; // @[IMemory.scala 502:50]
  assign _T_115 = io_aluop_i == 8'h44; // @[IMemory.scala 502:100]
  assign _T_116 = _T_114 | _T_115; // @[IMemory.scala 502:86]
  assign _T_117 = io_aluop_i == 8'h4c; // @[IMemory.scala 503:18]
  assign _T_118 = _T_116 | _T_117; // @[IMemory.scala 502:122]
  assign _T_119 = io_aluop_i == 8'h48; // @[IMemory.scala 503:54]
  assign _T_120 = _T_118 | _T_119; // @[IMemory.scala 503:40]
  assign _T_121 = io_aluop_i == 8'h70; // @[IMemory.scala 503:89]
  assign _T_122 = _T_120 | _T_121; // @[IMemory.scala 503:75]
  assign _T_123 = io_aluop_i == 8'h54; // @[IMemory.scala 504:18]
  assign _T_124 = _T_122 | _T_123; // @[IMemory.scala 503:111]
  assign _T_125 = io_aluop_i == 8'h79; // @[IMemory.scala 504:54]
  assign _T_126 = _T_124 | _T_125; // @[IMemory.scala 504:40]
  assign _T_127 = io_aluop_i == 8'h5c; // @[IMemory.scala 504:91]
  assign _T_128 = _T_126 | _T_127; // @[IMemory.scala 504:77]
  assign _T_129 = io_data_tlb_r_exception_i | io_data_tlb_w_exception_i; // @[IMemory.scala 506:38]
  assign _T_130 = io_cnt_i == 2'h0; // @[IMemory.scala 508:27]
  assign _T_135 = io_cnt_i == 2'h1; // @[IMemory.scala 530:27]
  assign _T_139 = io_original_data_i + io_reg2_i; // @[IMemory.scala 542:92]
  assign _T_141 = io_original_data_i ^ io_reg2_i; // @[IMemory.scala 543:92]
  assign _T_143 = io_original_data_i & io_reg2_i; // @[IMemory.scala 544:92]
  assign _T_145 = io_original_data_i | io_reg2_i; // @[IMemory.scala 545:92]
  assign _T_149 = $signed(io_original_data_i) < $signed(io_reg2_i); // @[IMemory.scala 546:103]
  assign _T_154 = $signed(io_original_data_i) > $signed(io_reg2_i); // @[IMemory.scala 547:103]
  assign _T_157 = io_original_data_i < io_reg2_i; // @[IMemory.scala 548:96]
  assign _T_160 = io_original_data_i > io_reg2_i; // @[IMemory.scala 549:96]
  assign _GEN_173 = _T_130 ? _T_4 : _T_135; // @[IMemory.scala 508:40]
  assign _GEN_176 = _T_130 ? 1'h0 : _T_135; // @[IMemory.scala 508:40]
  assign _GEN_177 = _T_130 | _T_135; // @[IMemory.scala 508:40]
  assign _GEN_180 = _T_130 & _T_4; // @[IMemory.scala 508:40]
  assign _GEN_188 = _T_129 ? 1'h0 : _GEN_173; // @[IMemory.scala 506:66]
  assign _GEN_191 = _T_129 ? 1'h0 : _GEN_176; // @[IMemory.scala 506:66]
  assign _GEN_192 = _T_129 ? 1'h0 : _GEN_177; // @[IMemory.scala 506:66]
  assign _GEN_195 = _T_129 ? 1'h0 : _GEN_180; // @[IMemory.scala 506:66]
  assign _GEN_203 = _T_128 & _GEN_188; // @[IMemory.scala 504:114]
  assign _GEN_206 = _T_128 & _GEN_191; // @[IMemory.scala 504:114]
  assign _GEN_207 = _T_128 & _GEN_192; // @[IMemory.scala 504:114]
  assign _GEN_210 = _T_128 & _GEN_195; // @[IMemory.scala 504:114]
  assign _GEN_312 = _T_81 & _GEN_21; // @[IMemory.scala 355:43]
  assign _GEN_479 = io_not_stall_i ? io_excepttype_i : 32'h0; // @[IMemory.scala 616:28]
  assign io_wd_o = io_rst_n ? wd_o : 5'h0; // @[IMemory.scala 116:11 IMemory.scala 590:11]
  assign io_wreg_o = io_rst_n ? wreg_o : 1'h0; // @[IMemory.scala 117:13 IMemory.scala 591:13]
  assign io_wdata_o = io_rst_n ? wdata_o : 32'h0; // @[IMemory.scala 118:14 IMemory.scala 592:14]
  assign io_LLbit_we_o = io_rst_n ? LLbit_we_o : 1'h0; // @[IMemory.scala 131:17 IMemory.scala 605:17]
  assign io_LLbit_value_o = io_rst_n ? LLbit_value_o : 1'h0; // @[IMemory.scala 133:20 IMemory.scala 607:20]
  assign io_LLbit_addr_o = io_rst_n ? LLbit_addr_o : 34'h0; // @[IMemory.scala 132:19 IMemory.scala 606:19]
  assign io_stallreq = io_stallreq_from_mem_i | stallreq_from_amo; // @[IMemory.scala 82:15 IMemory.scala 91:15]
  assign io_cnt_o = io_rst_n ? cnt_o : 2'h0; // @[IMemory.scala 135:12 IMemory.scala 609:12]
  assign io_original_data_o = io_rst_n ? original_data_o : 32'h0; // @[IMemory.scala 136:22 IMemory.scala 610:22]
  assign io_csr_reg_we_o = 1'h0; // @[IMemory.scala 120:19 IMemory.scala 594:19]
  assign io_csr_reg_addr_o = 12'h0; // @[IMemory.scala 121:21 IMemory.scala 595:21]
  assign io_csr_reg_data_o = 32'h0; // @[IMemory.scala 122:21 IMemory.scala 596:21]
  assign io_excepttype_o = io_rst_n ? _GEN_479 : 32'h0; // @[IMemory.scala 615:19 IMemory.scala 617:19 IMemory.scala 619:19]
  assign io_is_in_delayslot_o = io_is_in_delayslot_i; // @[IMemory.scala 79:24]
  assign io_current_inst_address_o = io_current_inst_address_i; // @[IMemory.scala 80:29]
  assign io_current_data_address_o = io_mem_addr_i; // @[IMemory.scala 81:29]
  assign io_not_stall_o = io_not_stall_i; // @[IMemory.scala 622:16]
  assign io_mem_addr_o = io_rst_n ? mem_addr_o : 32'h0; // @[IMemory.scala 124:17 IMemory.scala 598:17]
  assign io_mem_phy_addr_o = io_rst_n ? mem_phy_addr_o : 34'h0; // @[IMemory.scala 125:21 IMemory.scala 599:21]
  assign io_mem_we_o = io_rst_n ? mem_we_o : 1'h0; // @[IMemory.scala 126:15 IMemory.scala 600:15]
  assign io_mem_sel_o = io_rst_n ? mem_sel_o : 4'h0; // @[IMemory.scala 127:16 IMemory.scala 601:16]
  assign io_mem_data_o = io_rst_n ? mem_data_o : 32'h0; // @[IMemory.scala 128:17 IMemory.scala 541:66 IMemory.scala 550:40 IMemory.scala 602:17]
  assign io_mem_ce_o = io_rst_n ? mem_ce_o : 1'h0; // @[IMemory.scala 129:15 IMemory.scala 603:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stallreq_from_amo = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  wd_o = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  wreg_o = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  wdata_o = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mem_addr_o = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  mem_phy_addr_o = _RAND_5[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mem_we_o = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mem_sel_o = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_data_o = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  mem_ce_o = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  LLbit_we_o = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  LLbit_addr_o = _RAND_11[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  LLbit_value_o = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  cnt_o = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  original_data_o = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(*) begin
    if (~io_rst_n) begin
      stallreq_from_amo <= 1'h0;
    end else if (_T_2) begin
      stallreq_from_amo <= 1'h0;
    end else if (_T_31) begin
      stallreq_from_amo <= 1'h0;
    end else if (_T_52) begin
      stallreq_from_amo <= 1'h0;
    end else if (_T_67) begin
      stallreq_from_amo <= 1'h0;
    end else if (_T_78) begin
      stallreq_from_amo <= 1'h0;
    end else if (_T_81) begin
      stallreq_from_amo <= 1'h0;
    end else if (_T_84) begin
      stallreq_from_amo <= 1'h0;
    end else if (_T_96) begin
      stallreq_from_amo <= 1'h0;
    end else if (_T_103) begin
      stallreq_from_amo <= 1'h0;
    end else if (_T_106) begin
      stallreq_from_amo <= 1'h0;
    end else begin
      stallreq_from_amo <= _GEN_210;
    end
    if (~io_rst_n) begin
      wd_o <= 5'h0;
    end else if (~io_rst_n) begin
      wd_o <= 5'h0;
    end else begin
      wd_o <= io_wd_i;
    end
    if (~io_rst_n) begin
      wreg_o <= 1'h0;
    end else if (~io_rst_n) begin
      wreg_o <= 1'h0;
    end else begin
      wreg_o <= io_wreg_i;
    end
    if (~io_rst_n) begin
      wdata_o <= 32'h0;
    end else if (~io_rst_n) begin
      wdata_o <= 32'h0;
    end else if (_T_2) begin
      if (io_data_tlb_r_exception_i) begin
        wdata_o <= io_wdata_i;
      end else if (_T_4) begin
        wdata_o <= _T_9;
      end else if (_T_11) begin
        wdata_o <= _T_16;
      end else if (_T_18) begin
        wdata_o <= _T_23;
      end else if (_T_25) begin
        wdata_o <= _T_30;
      end else begin
        wdata_o <= 32'h0;
      end
    end else if (_T_31) begin
      if (io_data_tlb_r_exception_i) begin
        wdata_o <= io_wdata_i;
      end else if (_T_4) begin
        wdata_o <= _T_36;
      end else if (_T_11) begin
        wdata_o <= _T_41;
      end else if (_T_18) begin
        wdata_o <= _T_46;
      end else if (_T_25) begin
        wdata_o <= _T_51;
      end else begin
        wdata_o <= 32'h0;
      end
    end else if (_T_52) begin
      if (io_data_tlb_r_exception_i) begin
        wdata_o <= io_wdata_i;
      end else if (_T_4) begin
        wdata_o <= _T_59;
      end else if (_T_18) begin
        wdata_o <= _T_66;
      end else begin
        wdata_o <= 32'h0;
      end
    end else if (_T_67) begin
      if (io_data_tlb_r_exception_i) begin
        wdata_o <= io_wdata_i;
      end else if (_T_4) begin
        wdata_o <= _T_72;
      end else if (_T_18) begin
        wdata_o <= _T_77;
      end else begin
        wdata_o <= 32'h0;
      end
    end else if (_T_78) begin
      if (io_data_tlb_r_exception_i) begin
        wdata_o <= io_wdata_i;
      end else if (_T_4) begin
        wdata_o <= io_mem_data_i;
      end else begin
        wdata_o <= 32'h0;
      end
    end else if (_T_81) begin
      if (io_data_tlb_r_exception_i) begin
        wdata_o <= io_wdata_i;
      end else if (_T_4) begin
        wdata_o <= io_mem_data_i;
      end else begin
        wdata_o <= 32'h0;
      end
    end else if (_T_84) begin
      wdata_o <= io_wdata_i;
    end else if (_T_96) begin
      wdata_o <= io_wdata_i;
    end else if (_T_103) begin
      wdata_o <= io_wdata_i;
    end else if (_T_106) begin
      if (io_data_tlb_w_exception_i) begin
        wdata_o <= io_wdata_i;
      end else if (_T_109) begin
        wdata_o <= 32'h0;
      end else begin
        wdata_o <= 32'h1;
      end
    end else if (_T_128) begin
      if (_T_129) begin
        wdata_o <= io_wdata_i;
      end else if (_T_130) begin
        wdata_o <= io_wdata_i;
      end else if (_T_135) begin
        wdata_o <= io_original_data_i;
      end else begin
        wdata_o <= io_wdata_i;
      end
    end else begin
      wdata_o <= io_wdata_i;
    end
    if (~io_rst_n) begin
      mem_addr_o <= 32'h0;
    end else if (~io_rst_n) begin
      mem_addr_o <= 32'h0;
    end else if (_T_2) begin
      if (io_data_tlb_r_exception_i) begin
        mem_addr_o <= 32'h0;
      end else begin
        mem_addr_o <= io_mem_addr_i;
      end
    end else if (_T_31) begin
      if (io_data_tlb_r_exception_i) begin
        mem_addr_o <= 32'h0;
      end else begin
        mem_addr_o <= io_mem_addr_i;
      end
    end else if (_T_52) begin
      if (io_data_tlb_r_exception_i) begin
        mem_addr_o <= 32'h0;
      end else begin
        mem_addr_o <= io_mem_addr_i;
      end
    end else if (_T_67) begin
      if (io_data_tlb_r_exception_i) begin
        mem_addr_o <= 32'h0;
      end else begin
        mem_addr_o <= io_mem_addr_i;
      end
    end else if (_T_78) begin
      mem_addr_o <= _GEN_18;
    end else if (_T_81) begin
      mem_addr_o <= _GEN_18;
    end else if (_T_84) begin
      if (io_data_tlb_w_exception_i) begin
        mem_addr_o <= 32'h0;
      end else begin
        mem_addr_o <= io_mem_addr_i;
      end
    end else if (_T_96) begin
      if (io_data_tlb_w_exception_i) begin
        mem_addr_o <= 32'h0;
      end else begin
        mem_addr_o <= io_mem_addr_i;
      end
    end else if (_T_103) begin
      if (io_data_tlb_w_exception_i) begin
        mem_addr_o <= 32'h0;
      end else begin
        mem_addr_o <= io_mem_addr_i;
      end
    end else if (_T_106) begin
      if (io_data_tlb_w_exception_i) begin
        mem_addr_o <= 32'h0;
      end else begin
        mem_addr_o <= io_mem_addr_i;
      end
    end else if (_T_128) begin
      if (_T_129) begin
        mem_addr_o <= 32'h0;
      end else if (_T_130) begin
        mem_addr_o <= io_mem_addr_i;
      end else if (_T_135) begin
        mem_addr_o <= io_mem_addr_i;
      end else begin
        mem_addr_o <= 32'h0;
      end
    end else begin
      mem_addr_o <= 32'h0;
    end
    if (~io_rst_n) begin
      mem_phy_addr_o <= 34'h0;
    end else if (~io_rst_n) begin
      mem_phy_addr_o <= 34'h0;
    end else if (_T_2) begin
      if (io_data_tlb_r_exception_i) begin
        mem_phy_addr_o <= 34'h0;
      end else begin
        mem_phy_addr_o <= io_mem_phy_addr_i;
      end
    end else if (_T_31) begin
      if (io_data_tlb_r_exception_i) begin
        mem_phy_addr_o <= 34'h0;
      end else begin
        mem_phy_addr_o <= io_mem_phy_addr_i;
      end
    end else if (_T_52) begin
      if (io_data_tlb_r_exception_i) begin
        mem_phy_addr_o <= 34'h0;
      end else begin
        mem_phy_addr_o <= io_mem_phy_addr_i;
      end
    end else if (_T_67) begin
      if (io_data_tlb_r_exception_i) begin
        mem_phy_addr_o <= 34'h0;
      end else begin
        mem_phy_addr_o <= io_mem_phy_addr_i;
      end
    end else if (_T_78) begin
      mem_phy_addr_o <= _GEN_19;
    end else if (_T_81) begin
      mem_phy_addr_o <= _GEN_19;
    end else if (_T_84) begin
      if (io_data_tlb_w_exception_i) begin
        mem_phy_addr_o <= 34'h0;
      end else begin
        mem_phy_addr_o <= io_mem_phy_addr_i;
      end
    end else if (_T_96) begin
      if (io_data_tlb_w_exception_i) begin
        mem_phy_addr_o <= 34'h0;
      end else begin
        mem_phy_addr_o <= io_mem_phy_addr_i;
      end
    end else if (_T_103) begin
      if (io_data_tlb_w_exception_i) begin
        mem_phy_addr_o <= 34'h0;
      end else begin
        mem_phy_addr_o <= io_mem_phy_addr_i;
      end
    end else if (_T_106) begin
      if (io_data_tlb_w_exception_i) begin
        mem_phy_addr_o <= 34'h0;
      end else begin
        mem_phy_addr_o <= io_mem_phy_addr_i;
      end
    end else if (_T_128) begin
      if (_T_129) begin
        mem_phy_addr_o <= 34'h0;
      end else if (_T_130) begin
        mem_phy_addr_o <= io_mem_phy_addr_i;
      end else if (_T_135) begin
        mem_phy_addr_o <= io_mem_phy_addr_i;
      end else begin
        mem_phy_addr_o <= 34'h0;
      end
    end else begin
      mem_phy_addr_o <= 34'h0;
    end
    if (~io_rst_n) begin
      mem_we_o <= 1'h0;
    end else if (~io_rst_n) begin
      mem_we_o <= 1'h0;
    end else if (_T_2) begin
      mem_we_o <= 1'h0;
    end else if (_T_31) begin
      mem_we_o <= 1'h0;
    end else if (_T_52) begin
      mem_we_o <= 1'h0;
    end else if (_T_67) begin
      mem_we_o <= 1'h0;
    end else if (_T_78) begin
      mem_we_o <= 1'h0;
    end else if (_T_81) begin
      mem_we_o <= 1'h0;
    end else if (_T_84) begin
      if (io_data_tlb_w_exception_i) begin
        mem_we_o <= 1'h0;
      end else begin
        mem_we_o <= 1'h1;
      end
    end else if (_T_96) begin
      if (io_data_tlb_w_exception_i) begin
        mem_we_o <= 1'h0;
      end else begin
        mem_we_o <= 1'h1;
      end
    end else if (_T_103) begin
      if (io_data_tlb_w_exception_i) begin
        mem_we_o <= 1'h0;
      end else begin
        mem_we_o <= 1'h1;
      end
    end else if (_T_106) begin
      if (io_data_tlb_w_exception_i) begin
        mem_we_o <= 1'h0;
      end else begin
        mem_we_o <= 1'h1;
      end
    end else begin
      mem_we_o <= _GEN_206;
    end
    if (~io_rst_n) begin
      mem_sel_o <= 4'h0;
    end else if (~io_rst_n) begin
      mem_sel_o <= 4'h0;
    end else if (_T_2) begin
      if (io_data_tlb_r_exception_i) begin
        mem_sel_o <= 4'hf;
      end else if (_T_4) begin
        mem_sel_o <= 4'h1;
      end else if (_T_11) begin
        mem_sel_o <= 4'h2;
      end else if (_T_18) begin
        mem_sel_o <= 4'h4;
      end else if (_T_25) begin
        mem_sel_o <= 4'h8;
      end else begin
        mem_sel_o <= 4'h0;
      end
    end else if (_T_31) begin
      if (io_data_tlb_r_exception_i) begin
        mem_sel_o <= 4'hf;
      end else if (_T_4) begin
        mem_sel_o <= 4'h1;
      end else if (_T_11) begin
        mem_sel_o <= 4'h2;
      end else if (_T_18) begin
        mem_sel_o <= 4'h4;
      end else if (_T_25) begin
        mem_sel_o <= 4'h8;
      end else begin
        mem_sel_o <= 4'h0;
      end
    end else if (_T_52) begin
      if (io_data_tlb_r_exception_i) begin
        mem_sel_o <= 4'hf;
      end else if (_T_4) begin
        mem_sel_o <= 4'h3;
      end else if (_T_18) begin
        mem_sel_o <= 4'hc;
      end else begin
        mem_sel_o <= 4'h0;
      end
    end else if (_T_67) begin
      if (io_data_tlb_r_exception_i) begin
        mem_sel_o <= 4'hf;
      end else if (_T_4) begin
        mem_sel_o <= 4'h3;
      end else if (_T_18) begin
        mem_sel_o <= 4'hc;
      end else begin
        mem_sel_o <= 4'h0;
      end
    end else if (_T_78) begin
      if (io_data_tlb_r_exception_i) begin
        mem_sel_o <= 4'hf;
      end else if (_T_4) begin
        mem_sel_o <= 4'hf;
      end else begin
        mem_sel_o <= 4'h0;
      end
    end else if (_T_81) begin
      if (io_data_tlb_r_exception_i) begin
        mem_sel_o <= 4'hf;
      end else if (_T_4) begin
        mem_sel_o <= 4'hf;
      end else begin
        mem_sel_o <= 4'h0;
      end
    end else if (_T_84) begin
      if (io_data_tlb_w_exception_i) begin
        mem_sel_o <= 4'hf;
      end else if (_T_4) begin
        mem_sel_o <= 4'h1;
      end else if (_T_11) begin
        mem_sel_o <= 4'h2;
      end else if (_T_18) begin
        mem_sel_o <= 4'h4;
      end else if (_T_25) begin
        mem_sel_o <= 4'h8;
      end else begin
        mem_sel_o <= 4'h0;
      end
    end else if (_T_96) begin
      if (io_data_tlb_w_exception_i) begin
        mem_sel_o <= 4'hf;
      end else if (_T_4) begin
        mem_sel_o <= 4'h3;
      end else if (_T_18) begin
        mem_sel_o <= 4'hc;
      end else begin
        mem_sel_o <= 4'h0;
      end
    end else if (_T_103) begin
      if (io_data_tlb_w_exception_i) begin
        mem_sel_o <= 4'hf;
      end else if (_T_4) begin
        mem_sel_o <= 4'hf;
      end else begin
        mem_sel_o <= 4'h0;
      end
    end else if (_T_106) begin
      if (io_data_tlb_w_exception_i) begin
        mem_sel_o <= 4'hf;
      end else if (_T_109) begin
        if (_T_4) begin
          mem_sel_o <= 4'hf;
        end else begin
          mem_sel_o <= 4'h0;
        end
      end else begin
        mem_sel_o <= 4'hf;
      end
    end else if (_T_128) begin
      if (_T_129) begin
        mem_sel_o <= 4'hf;
      end else if (_T_130) begin
        mem_sel_o <= _GEN_70;
      end else begin
        mem_sel_o <= 4'hf;
      end
    end else begin
      mem_sel_o <= 4'hf;
    end
    if (~io_rst_n) begin
      mem_data_o <= 32'h0;
    end else if (~io_rst_n) begin
      mem_data_o <= 32'h0;
    end else if (_T_2) begin
      mem_data_o <= 32'h0;
    end else if (_T_31) begin
      mem_data_o <= 32'h0;
    end else if (_T_52) begin
      mem_data_o <= 32'h0;
    end else if (_T_67) begin
      mem_data_o <= 32'h0;
    end else if (_T_78) begin
      mem_data_o <= 32'h0;
    end else if (_T_81) begin
      mem_data_o <= 32'h0;
    end else if (_T_84) begin
      if (io_data_tlb_w_exception_i) begin
        mem_data_o <= 32'h0;
      end else begin
        mem_data_o <= _T_87;
      end
    end else if (_T_96) begin
      if (io_data_tlb_w_exception_i) begin
        mem_data_o <= 32'h0;
      end else begin
        mem_data_o <= _T_98;
      end
    end else if (_T_103) begin
      if (io_data_tlb_w_exception_i) begin
        mem_data_o <= 32'h0;
      end else begin
        mem_data_o <= io_reg2_i;
      end
    end else if (_T_106) begin
      if (io_data_tlb_w_exception_i) begin
        mem_data_o <= 32'h0;
      end else if (_T_109) begin
        mem_data_o <= io_reg2_i;
      end else begin
        mem_data_o <= 32'h0;
      end
    end else if (_T_128) begin
      if (_T_129) begin
        mem_data_o <= 32'h0;
      end else if (_T_130) begin
        mem_data_o <= 32'h0;
      end else if (_T_135) begin
        if (_T_112) begin
          mem_data_o <= 32'h0;
        end else if (_T_113) begin
          mem_data_o <= _T_139;
        end else if (_T_115) begin
          mem_data_o <= _T_141;
        end else if (_T_117) begin
          mem_data_o <= _T_143;
        end else if (_T_119) begin
          mem_data_o <= _T_145;
        end else if (_T_121) begin
          if (_T_149) begin
            mem_data_o <= io_original_data_i;
          end else begin
            mem_data_o <= io_reg2_i;
          end
        end else if (_T_123) begin
          if (_T_154) begin
            mem_data_o <= io_original_data_i;
          end else begin
            mem_data_o <= io_reg2_i;
          end
        end else if (_T_125) begin
          if (_T_157) begin
            mem_data_o <= io_original_data_i;
          end else begin
            mem_data_o <= io_reg2_i;
          end
        end else if (_T_127) begin
          if (_T_160) begin
            mem_data_o <= io_original_data_i;
          end else begin
            mem_data_o <= io_reg2_i;
          end
        end else begin
          mem_data_o <= 32'h0;
        end
      end else begin
        mem_data_o <= 32'h0;
      end
    end else begin
      mem_data_o <= 32'h0;
    end
    if (~io_rst_n) begin
      mem_ce_o <= 1'h0;
    end else if (~io_rst_n) begin
      mem_ce_o <= 1'h0;
    end else if (_T_2) begin
      if (io_data_tlb_r_exception_i) begin
        mem_ce_o <= 1'h0;
      end else begin
        mem_ce_o <= _GEN_14;
      end
    end else if (_T_31) begin
      if (io_data_tlb_r_exception_i) begin
        mem_ce_o <= 1'h0;
      end else begin
        mem_ce_o <= _GEN_14;
      end
    end else if (_T_52) begin
      if (io_data_tlb_r_exception_i) begin
        mem_ce_o <= 1'h0;
      end else begin
        mem_ce_o <= _GEN_51;
      end
    end else if (_T_67) begin
      if (io_data_tlb_r_exception_i) begin
        mem_ce_o <= 1'h0;
      end else begin
        mem_ce_o <= _GEN_51;
      end
    end else if (_T_78) begin
      if (io_data_tlb_r_exception_i) begin
        mem_ce_o <= 1'h0;
      end else begin
        mem_ce_o <= _T_4;
      end
    end else if (_T_81) begin
      if (io_data_tlb_r_exception_i) begin
        mem_ce_o <= 1'h0;
      end else begin
        mem_ce_o <= _T_4;
      end
    end else if (_T_84) begin
      if (io_data_tlb_w_exception_i) begin
        mem_ce_o <= 1'h0;
      end else begin
        mem_ce_o <= _GEN_14;
      end
    end else if (_T_96) begin
      if (io_data_tlb_w_exception_i) begin
        mem_ce_o <= 1'h0;
      end else begin
        mem_ce_o <= _GEN_51;
      end
    end else if (_T_103) begin
      if (io_data_tlb_w_exception_i) begin
        mem_ce_o <= 1'h0;
      end else begin
        mem_ce_o <= _T_4;
      end
    end else if (_T_106) begin
      if (io_data_tlb_w_exception_i) begin
        mem_ce_o <= 1'h0;
      end else begin
        mem_ce_o <= _GEN_124;
      end
    end else begin
      mem_ce_o <= _GEN_203;
    end
    if (~io_rst_n) begin
      LLbit_we_o <= 1'h0;
    end else if (~io_rst_n) begin
      LLbit_we_o <= 1'h0;
    end else if (_T_2) begin
      if (io_data_tlb_r_exception_i) begin
        LLbit_we_o <= 1'h0;
      end else begin
        LLbit_we_o <= 1'h1;
      end
    end else if (_T_31) begin
      if (io_data_tlb_r_exception_i) begin
        LLbit_we_o <= 1'h0;
      end else begin
        LLbit_we_o <= 1'h1;
      end
    end else if (_T_52) begin
      if (io_data_tlb_r_exception_i) begin
        LLbit_we_o <= 1'h0;
      end else begin
        LLbit_we_o <= 1'h1;
      end
    end else if (_T_67) begin
      if (io_data_tlb_r_exception_i) begin
        LLbit_we_o <= 1'h0;
      end else begin
        LLbit_we_o <= 1'h1;
      end
    end else if (_T_78) begin
      LLbit_we_o <= _GEN_21;
    end else if (_T_81) begin
      LLbit_we_o <= _GEN_21;
    end else if (_T_84) begin
      LLbit_we_o <= _GEN_101;
    end else if (_T_96) begin
      LLbit_we_o <= _GEN_101;
    end else if (_T_103) begin
      LLbit_we_o <= _GEN_101;
    end else if (_T_106) begin
      LLbit_we_o <= _GEN_101;
    end else begin
      LLbit_we_o <= _GEN_207;
    end
    if (~io_rst_n) begin
      LLbit_addr_o <= 34'h0;
    end else if (~io_rst_n) begin
      LLbit_addr_o <= 34'h0;
    end else if (_T_2) begin
      LLbit_addr_o <= 34'h0;
    end else if (_T_31) begin
      LLbit_addr_o <= 34'h0;
    end else if (_T_52) begin
      LLbit_addr_o <= 34'h0;
    end else if (_T_67) begin
      LLbit_addr_o <= 34'h0;
    end else if (_T_78) begin
      LLbit_addr_o <= 34'h0;
    end else if (_T_81) begin
      LLbit_addr_o <= _GEN_19;
    end else begin
      LLbit_addr_o <= 34'h0;
    end
    if (~io_rst_n) begin
      LLbit_value_o <= 1'h0;
    end else if (~io_rst_n) begin
      LLbit_value_o <= 1'h0;
    end else if (_T_2) begin
      LLbit_value_o <= 1'h0;
    end else if (_T_31) begin
      LLbit_value_o <= 1'h0;
    end else if (_T_52) begin
      LLbit_value_o <= 1'h0;
    end else if (_T_67) begin
      LLbit_value_o <= 1'h0;
    end else if (_T_78) begin
      LLbit_value_o <= 1'h0;
    end else begin
      LLbit_value_o <= _GEN_312;
    end
    if (~io_rst_n) begin
      cnt_o <= 2'h0;
    end else if (~io_rst_n) begin
      cnt_o <= 2'h0;
    end else if (_T_2) begin
      cnt_o <= 2'h0;
    end else if (_T_31) begin
      cnt_o <= 2'h0;
    end else if (_T_52) begin
      cnt_o <= 2'h0;
    end else if (_T_67) begin
      cnt_o <= 2'h0;
    end else if (_T_78) begin
      cnt_o <= 2'h0;
    end else if (_T_81) begin
      cnt_o <= 2'h0;
    end else if (_T_84) begin
      cnt_o <= 2'h0;
    end else if (_T_96) begin
      cnt_o <= 2'h0;
    end else if (_T_103) begin
      cnt_o <= 2'h0;
    end else if (_T_106) begin
      cnt_o <= 2'h0;
    end else if (_T_128) begin
      if (_T_129) begin
        cnt_o <= 2'h0;
      end else if (_T_130) begin
        if (io_stallreq_from_mem_i) begin
          cnt_o <= 2'h0;
        end else begin
          cnt_o <= 2'h1;
        end
      end else if (_T_135) begin
        cnt_o <= 2'h1;
      end else begin
        cnt_o <= 2'h0;
      end
    end else begin
      cnt_o <= 2'h0;
    end
    if (~io_rst_n) begin
      original_data_o <= 32'h0;
    end else if (~io_rst_n) begin
      original_data_o <= 32'h0;
    end else if (_T_2) begin
      original_data_o <= 32'h0;
    end else if (_T_31) begin
      original_data_o <= 32'h0;
    end else if (_T_52) begin
      original_data_o <= 32'h0;
    end else if (_T_67) begin
      original_data_o <= 32'h0;
    end else if (_T_78) begin
      original_data_o <= 32'h0;
    end else if (_T_81) begin
      original_data_o <= 32'h0;
    end else if (_T_84) begin
      original_data_o <= 32'h0;
    end else if (_T_96) begin
      original_data_o <= 32'h0;
    end else if (_T_103) begin
      original_data_o <= 32'h0;
    end else if (_T_106) begin
      original_data_o <= 32'h0;
    end else if (_T_128) begin
      if (_T_129) begin
        original_data_o <= 32'h0;
      end else if (_T_130) begin
        original_data_o <= io_mem_data_i;
      end else if (_T_135) begin
        original_data_o <= io_original_data_i;
      end else begin
        original_data_o <= 32'h0;
      end
    end else begin
      original_data_o <= 32'h0;
    end
  end
endmodule
