module mmu_conv_chisel(
  input         io_rst_n,
  input  [31:0] io_tlb0_vpn_i,
  input  [31:0] io_tlb0_mask_i,
  input  [31:0] io_tlb0_pte_i,
  input  [31:0] io_tlb1_vpn_i,
  input  [31:0] io_tlb1_mask_i,
  input  [31:0] io_tlb1_pte_i,
  input  [31:0] io_tlb2_vpn_i,
  input  [31:0] io_tlb2_mask_i,
  input  [31:0] io_tlb2_pte_i,
  input  [31:0] io_tlb3_vpn_i,
  input  [31:0] io_tlb3_mask_i,
  input  [31:0] io_tlb3_pte_i,
  input  [31:0] io_tlb4_vpn_i,
  input  [31:0] io_tlb4_mask_i,
  input  [31:0] io_tlb4_pte_i,
  input  [31:0] io_tlb5_vpn_i,
  input  [31:0] io_tlb5_mask_i,
  input  [31:0] io_tlb5_pte_i,
  input  [31:0] io_tlb6_vpn_i,
  input  [31:0] io_tlb6_mask_i,
  input  [31:0] io_tlb6_pte_i,
  input  [31:0] io_tlb7_vpn_i,
  input  [31:0] io_tlb7_mask_i,
  input  [31:0] io_tlb7_pte_i,
  input  [31:0] io_tlb8_vpn_i,
  input  [31:0] io_tlb8_mask_i,
  input  [31:0] io_tlb8_pte_i,
  input  [31:0] io_tlb9_vpn_i,
  input  [31:0] io_tlb9_mask_i,
  input  [31:0] io_tlb9_pte_i,
  input  [31:0] io_tlb10_vpn_i,
  input  [31:0] io_tlb10_mask_i,
  input  [31:0] io_tlb10_pte_i,
  input  [31:0] io_tlb11_vpn_i,
  input  [31:0] io_tlb11_mask_i,
  input  [31:0] io_tlb11_pte_i,
  input  [31:0] io_tlb12_vpn_i,
  input  [31:0] io_tlb12_mask_i,
  input  [31:0] io_tlb12_pte_i,
  input  [31:0] io_tlb13_vpn_i,
  input  [31:0] io_tlb13_mask_i,
  input  [31:0] io_tlb13_pte_i,
  input  [31:0] io_tlb14_vpn_i,
  input  [31:0] io_tlb14_mask_i,
  input  [31:0] io_tlb14_pte_i,
  input  [31:0] io_tlb15_vpn_i,
  input  [31:0] io_tlb15_mask_i,
  input  [31:0] io_tlb15_pte_i,
  input  [4:0]  io_vm_i,
  input  [1:0]  io_prv_i,
  input         io_mxr_i,
  input         io_ce_i,
  input         io_ex_i,
  input         io_we_i,
  input  [31:0] io_vir_addr_i,
  output [33:0] io_phy_addr_o,
  output        io_tlb_exception_o,
  output        io_tlb_update_o,
  output [3:0]  io_hit_index_o
);
  reg [31:0] tlb_vpn_0; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_0;
  reg [31:0] tlb_vpn_1; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_1;
  reg [31:0] tlb_vpn_2; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_2;
  reg [31:0] tlb_vpn_3; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_3;
  reg [31:0] tlb_vpn_4; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_4;
  reg [31:0] tlb_vpn_5; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_5;
  reg [31:0] tlb_vpn_6; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_6;
  reg [31:0] tlb_vpn_7; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_7;
  reg [31:0] tlb_vpn_8; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_8;
  reg [31:0] tlb_vpn_9; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_9;
  reg [31:0] tlb_vpn_10; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_10;
  reg [31:0] tlb_vpn_11; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_11;
  reg [31:0] tlb_vpn_12; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_12;
  reg [31:0] tlb_vpn_13; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_13;
  reg [31:0] tlb_vpn_14; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_14;
  reg [31:0] tlb_vpn_15; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_15;
  reg [31:0] tlb_pte_0; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_16;
  reg [31:0] tlb_pte_1; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_17;
  reg [31:0] tlb_pte_2; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_18;
  reg [31:0] tlb_pte_3; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_19;
  reg [31:0] tlb_pte_4; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_20;
  reg [31:0] tlb_pte_5; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_21;
  reg [31:0] tlb_pte_6; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_22;
  reg [31:0] tlb_pte_7; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_23;
  reg [31:0] tlb_pte_8; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_24;
  reg [31:0] tlb_pte_9; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_25;
  reg [31:0] tlb_pte_10; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_26;
  reg [31:0] tlb_pte_11; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_27;
  reg [31:0] tlb_pte_12; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_28;
  reg [31:0] tlb_pte_13; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_29;
  reg [31:0] tlb_pte_14; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_30;
  reg [31:0] tlb_pte_15; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_31;
  reg [31:0] tlb_mask_0; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_32;
  reg [31:0] tlb_mask_1; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_33;
  reg [31:0] tlb_mask_2; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_34;
  reg [31:0] tlb_mask_3; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_35;
  reg [31:0] tlb_mask_4; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_36;
  reg [31:0] tlb_mask_5; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_37;
  reg [31:0] tlb_mask_6; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_38;
  reg [31:0] tlb_mask_7; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_39;
  reg [31:0] tlb_mask_8; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_40;
  reg [31:0] tlb_mask_9; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_41;
  reg [31:0] tlb_mask_10; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_42;
  reg [31:0] tlb_mask_11; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_43;
  reg [31:0] tlb_mask_12; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_44;
  reg [31:0] tlb_mask_13; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_45;
  reg [31:0] tlb_mask_14; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_46;
  reg [31:0] tlb_mask_15; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_47;
  reg [33:0] phy_addr_0; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_48;
  reg [33:0] phy_addr_1; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_49;
  reg [33:0] phy_addr_2; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_50;
  reg [33:0] phy_addr_3; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_51;
  reg [33:0] phy_addr_4; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_52;
  reg [33:0] phy_addr_5; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_53;
  reg [33:0] phy_addr_6; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_54;
  reg [33:0] phy_addr_7; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_55;
  reg [33:0] phy_addr_8; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_56;
  reg [33:0] phy_addr_9; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_57;
  reg [33:0] phy_addr_10; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_58;
  reg [33:0] phy_addr_11; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_59;
  reg [33:0] phy_addr_12; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_60;
  reg [33:0] phy_addr_13; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_61;
  reg [33:0] phy_addr_14; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_62;
  reg [33:0] phy_addr_15; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_63;
  wire  _T; // @[mmu_conv.scala 109:18]
  wire  _T_1; // @[mmu_conv.scala 112:24]
  wire [31:0] _T_2; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_3; // @[mmu_conv.scala 113:64]
  wire  _T_4; // @[mmu_conv.scala 113:48]
  wire  _GEN_0; // @[mmu_conv.scala 112:50]
  wire  _GEN_1; // @[mmu_conv.scala 109:45]
  wire  hit_0; // @[mmu_conv.scala 119:32]
  wire  _GEN_3; // @[mmu_conv.scala 126:35]
  wire  _GEN_4; // @[mmu_conv.scala 129:35]
  wire  _GEN_5; // @[mmu_conv.scala 130:35]
  wire  _T_19; // @[mmu_conv.scala 134:36]
  wire  _GEN_6; // @[mmu_conv.scala 134:61]
  wire  _GEN_7; // @[mmu_conv.scala 138:36]
  wire  _GEN_8; // @[mmu_conv.scala 133:21]
  wire  _GEN_9; // @[mmu_conv.scala 128:42]
  wire  protect_exception_0; // @[mmu_conv.scala 125:18]
  wire  _GEN_11; // @[mmu_conv.scala 145:32]
  wire  _T_28; // @[mmu_conv.scala 148:36]
  wire  update_exception_0; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_29; // @[Cat.scala 29:58]
  wire [33:0] _GEN_286; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_30; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_32; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_287; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_36; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_37; // @[mmu_conv.scala 113:64]
  wire  _T_38; // @[mmu_conv.scala 113:48]
  wire  _GEN_13; // @[mmu_conv.scala 112:50]
  wire  _GEN_14; // @[mmu_conv.scala 109:45]
  wire  hit_1; // @[mmu_conv.scala 119:32]
  wire  _GEN_16; // @[mmu_conv.scala 126:35]
  wire  _GEN_17; // @[mmu_conv.scala 129:35]
  wire  _GEN_18; // @[mmu_conv.scala 130:35]
  wire  _T_53; // @[mmu_conv.scala 134:36]
  wire  _GEN_19; // @[mmu_conv.scala 134:61]
  wire  _GEN_20; // @[mmu_conv.scala 138:36]
  wire  _GEN_21; // @[mmu_conv.scala 133:21]
  wire  _GEN_22; // @[mmu_conv.scala 128:42]
  wire  protect_exception_1; // @[mmu_conv.scala 125:18]
  wire  _GEN_24; // @[mmu_conv.scala 145:32]
  wire  _T_62; // @[mmu_conv.scala 148:36]
  wire  update_exception_1; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_63; // @[Cat.scala 29:58]
  wire [33:0] _GEN_288; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_64; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_66; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_289; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_70; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_71; // @[mmu_conv.scala 113:64]
  wire  _T_72; // @[mmu_conv.scala 113:48]
  wire  _GEN_26; // @[mmu_conv.scala 112:50]
  wire  _GEN_27; // @[mmu_conv.scala 109:45]
  wire  hit_2; // @[mmu_conv.scala 119:32]
  wire  _GEN_29; // @[mmu_conv.scala 126:35]
  wire  _GEN_30; // @[mmu_conv.scala 129:35]
  wire  _GEN_31; // @[mmu_conv.scala 130:35]
  wire  _T_87; // @[mmu_conv.scala 134:36]
  wire  _GEN_32; // @[mmu_conv.scala 134:61]
  wire  _GEN_33; // @[mmu_conv.scala 138:36]
  wire  _GEN_34; // @[mmu_conv.scala 133:21]
  wire  _GEN_35; // @[mmu_conv.scala 128:42]
  wire  protect_exception_2; // @[mmu_conv.scala 125:18]
  wire  _GEN_37; // @[mmu_conv.scala 145:32]
  wire  _T_96; // @[mmu_conv.scala 148:36]
  wire  update_exception_2; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_97; // @[Cat.scala 29:58]
  wire [33:0] _GEN_290; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_98; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_100; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_291; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_104; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_105; // @[mmu_conv.scala 113:64]
  wire  _T_106; // @[mmu_conv.scala 113:48]
  wire  _GEN_39; // @[mmu_conv.scala 112:50]
  wire  _GEN_40; // @[mmu_conv.scala 109:45]
  wire  hit_3; // @[mmu_conv.scala 119:32]
  wire  _GEN_42; // @[mmu_conv.scala 126:35]
  wire  _GEN_43; // @[mmu_conv.scala 129:35]
  wire  _GEN_44; // @[mmu_conv.scala 130:35]
  wire  _T_121; // @[mmu_conv.scala 134:36]
  wire  _GEN_45; // @[mmu_conv.scala 134:61]
  wire  _GEN_46; // @[mmu_conv.scala 138:36]
  wire  _GEN_47; // @[mmu_conv.scala 133:21]
  wire  _GEN_48; // @[mmu_conv.scala 128:42]
  wire  protect_exception_3; // @[mmu_conv.scala 125:18]
  wire  _GEN_50; // @[mmu_conv.scala 145:32]
  wire  _T_130; // @[mmu_conv.scala 148:36]
  wire  update_exception_3; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_131; // @[Cat.scala 29:58]
  wire [33:0] _GEN_292; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_132; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_134; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_293; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_138; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_139; // @[mmu_conv.scala 113:64]
  wire  _T_140; // @[mmu_conv.scala 113:48]
  wire  _GEN_52; // @[mmu_conv.scala 112:50]
  wire  _GEN_53; // @[mmu_conv.scala 109:45]
  wire  hit_4; // @[mmu_conv.scala 119:32]
  wire  _GEN_55; // @[mmu_conv.scala 126:35]
  wire  _GEN_56; // @[mmu_conv.scala 129:35]
  wire  _GEN_57; // @[mmu_conv.scala 130:35]
  wire  _T_155; // @[mmu_conv.scala 134:36]
  wire  _GEN_58; // @[mmu_conv.scala 134:61]
  wire  _GEN_59; // @[mmu_conv.scala 138:36]
  wire  _GEN_60; // @[mmu_conv.scala 133:21]
  wire  _GEN_61; // @[mmu_conv.scala 128:42]
  wire  protect_exception_4; // @[mmu_conv.scala 125:18]
  wire  _GEN_63; // @[mmu_conv.scala 145:32]
  wire  _T_164; // @[mmu_conv.scala 148:36]
  wire  update_exception_4; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_165; // @[Cat.scala 29:58]
  wire [33:0] _GEN_294; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_166; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_168; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_295; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_172; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_173; // @[mmu_conv.scala 113:64]
  wire  _T_174; // @[mmu_conv.scala 113:48]
  wire  _GEN_65; // @[mmu_conv.scala 112:50]
  wire  _GEN_66; // @[mmu_conv.scala 109:45]
  wire  hit_5; // @[mmu_conv.scala 119:32]
  wire  _GEN_68; // @[mmu_conv.scala 126:35]
  wire  _GEN_69; // @[mmu_conv.scala 129:35]
  wire  _GEN_70; // @[mmu_conv.scala 130:35]
  wire  _T_189; // @[mmu_conv.scala 134:36]
  wire  _GEN_71; // @[mmu_conv.scala 134:61]
  wire  _GEN_72; // @[mmu_conv.scala 138:36]
  wire  _GEN_73; // @[mmu_conv.scala 133:21]
  wire  _GEN_74; // @[mmu_conv.scala 128:42]
  wire  protect_exception_5; // @[mmu_conv.scala 125:18]
  wire  _GEN_76; // @[mmu_conv.scala 145:32]
  wire  _T_198; // @[mmu_conv.scala 148:36]
  wire  update_exception_5; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_199; // @[Cat.scala 29:58]
  wire [33:0] _GEN_296; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_200; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_202; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_297; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_206; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_207; // @[mmu_conv.scala 113:64]
  wire  _T_208; // @[mmu_conv.scala 113:48]
  wire  _GEN_78; // @[mmu_conv.scala 112:50]
  wire  _GEN_79; // @[mmu_conv.scala 109:45]
  wire  hit_6; // @[mmu_conv.scala 119:32]
  wire  _GEN_81; // @[mmu_conv.scala 126:35]
  wire  _GEN_82; // @[mmu_conv.scala 129:35]
  wire  _GEN_83; // @[mmu_conv.scala 130:35]
  wire  _T_223; // @[mmu_conv.scala 134:36]
  wire  _GEN_84; // @[mmu_conv.scala 134:61]
  wire  _GEN_85; // @[mmu_conv.scala 138:36]
  wire  _GEN_86; // @[mmu_conv.scala 133:21]
  wire  _GEN_87; // @[mmu_conv.scala 128:42]
  wire  protect_exception_6; // @[mmu_conv.scala 125:18]
  wire  _GEN_89; // @[mmu_conv.scala 145:32]
  wire  _T_232; // @[mmu_conv.scala 148:36]
  wire  update_exception_6; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_233; // @[Cat.scala 29:58]
  wire [33:0] _GEN_298; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_234; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_236; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_299; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_240; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_241; // @[mmu_conv.scala 113:64]
  wire  _T_242; // @[mmu_conv.scala 113:48]
  wire  _GEN_91; // @[mmu_conv.scala 112:50]
  wire  _GEN_92; // @[mmu_conv.scala 109:45]
  wire  hit_7; // @[mmu_conv.scala 119:32]
  wire  _GEN_94; // @[mmu_conv.scala 126:35]
  wire  _GEN_95; // @[mmu_conv.scala 129:35]
  wire  _GEN_96; // @[mmu_conv.scala 130:35]
  wire  _T_257; // @[mmu_conv.scala 134:36]
  wire  _GEN_97; // @[mmu_conv.scala 134:61]
  wire  _GEN_98; // @[mmu_conv.scala 138:36]
  wire  _GEN_99; // @[mmu_conv.scala 133:21]
  wire  _GEN_100; // @[mmu_conv.scala 128:42]
  wire  protect_exception_7; // @[mmu_conv.scala 125:18]
  wire  _GEN_102; // @[mmu_conv.scala 145:32]
  wire  _T_266; // @[mmu_conv.scala 148:36]
  wire  update_exception_7; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_267; // @[Cat.scala 29:58]
  wire [33:0] _GEN_300; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_268; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_270; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_301; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_274; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_275; // @[mmu_conv.scala 113:64]
  wire  _T_276; // @[mmu_conv.scala 113:48]
  wire  _GEN_104; // @[mmu_conv.scala 112:50]
  wire  _GEN_105; // @[mmu_conv.scala 109:45]
  wire  hit_8; // @[mmu_conv.scala 119:32]
  wire  _GEN_107; // @[mmu_conv.scala 126:35]
  wire  _GEN_108; // @[mmu_conv.scala 129:35]
  wire  _GEN_109; // @[mmu_conv.scala 130:35]
  wire  _T_291; // @[mmu_conv.scala 134:36]
  wire  _GEN_110; // @[mmu_conv.scala 134:61]
  wire  _GEN_111; // @[mmu_conv.scala 138:36]
  wire  _GEN_112; // @[mmu_conv.scala 133:21]
  wire  _GEN_113; // @[mmu_conv.scala 128:42]
  wire  protect_exception_8; // @[mmu_conv.scala 125:18]
  wire  _GEN_115; // @[mmu_conv.scala 145:32]
  wire  _T_300; // @[mmu_conv.scala 148:36]
  wire  update_exception_8; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_301; // @[Cat.scala 29:58]
  wire [33:0] _GEN_302; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_302; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_304; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_303; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_308; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_309; // @[mmu_conv.scala 113:64]
  wire  _T_310; // @[mmu_conv.scala 113:48]
  wire  _GEN_117; // @[mmu_conv.scala 112:50]
  wire  _GEN_118; // @[mmu_conv.scala 109:45]
  wire  hit_9; // @[mmu_conv.scala 119:32]
  wire  _GEN_120; // @[mmu_conv.scala 126:35]
  wire  _GEN_121; // @[mmu_conv.scala 129:35]
  wire  _GEN_122; // @[mmu_conv.scala 130:35]
  wire  _T_325; // @[mmu_conv.scala 134:36]
  wire  _GEN_123; // @[mmu_conv.scala 134:61]
  wire  _GEN_124; // @[mmu_conv.scala 138:36]
  wire  _GEN_125; // @[mmu_conv.scala 133:21]
  wire  _GEN_126; // @[mmu_conv.scala 128:42]
  wire  protect_exception_9; // @[mmu_conv.scala 125:18]
  wire  _GEN_128; // @[mmu_conv.scala 145:32]
  wire  _T_334; // @[mmu_conv.scala 148:36]
  wire  update_exception_9; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_335; // @[Cat.scala 29:58]
  wire [33:0] _GEN_304; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_336; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_338; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_305; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_342; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_343; // @[mmu_conv.scala 113:64]
  wire  _T_344; // @[mmu_conv.scala 113:48]
  wire  _GEN_130; // @[mmu_conv.scala 112:50]
  wire  _GEN_131; // @[mmu_conv.scala 109:45]
  wire  hit_10; // @[mmu_conv.scala 119:32]
  wire  _GEN_133; // @[mmu_conv.scala 126:35]
  wire  _GEN_134; // @[mmu_conv.scala 129:35]
  wire  _GEN_135; // @[mmu_conv.scala 130:35]
  wire  _T_359; // @[mmu_conv.scala 134:36]
  wire  _GEN_136; // @[mmu_conv.scala 134:61]
  wire  _GEN_137; // @[mmu_conv.scala 138:36]
  wire  _GEN_138; // @[mmu_conv.scala 133:21]
  wire  _GEN_139; // @[mmu_conv.scala 128:42]
  wire  protect_exception_10; // @[mmu_conv.scala 125:18]
  wire  _GEN_141; // @[mmu_conv.scala 145:32]
  wire  _T_368; // @[mmu_conv.scala 148:36]
  wire  update_exception_10; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_369; // @[Cat.scala 29:58]
  wire [33:0] _GEN_306; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_370; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_372; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_307; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_376; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_377; // @[mmu_conv.scala 113:64]
  wire  _T_378; // @[mmu_conv.scala 113:48]
  wire  _GEN_143; // @[mmu_conv.scala 112:50]
  wire  _GEN_144; // @[mmu_conv.scala 109:45]
  wire  hit_11; // @[mmu_conv.scala 119:32]
  wire  _GEN_146; // @[mmu_conv.scala 126:35]
  wire  _GEN_147; // @[mmu_conv.scala 129:35]
  wire  _GEN_148; // @[mmu_conv.scala 130:35]
  wire  _T_393; // @[mmu_conv.scala 134:36]
  wire  _GEN_149; // @[mmu_conv.scala 134:61]
  wire  _GEN_150; // @[mmu_conv.scala 138:36]
  wire  _GEN_151; // @[mmu_conv.scala 133:21]
  wire  _GEN_152; // @[mmu_conv.scala 128:42]
  wire  protect_exception_11; // @[mmu_conv.scala 125:18]
  wire  _GEN_154; // @[mmu_conv.scala 145:32]
  wire  _T_402; // @[mmu_conv.scala 148:36]
  wire  update_exception_11; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_403; // @[Cat.scala 29:58]
  wire [33:0] _GEN_308; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_404; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_406; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_309; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_410; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_411; // @[mmu_conv.scala 113:64]
  wire  _T_412; // @[mmu_conv.scala 113:48]
  wire  _GEN_156; // @[mmu_conv.scala 112:50]
  wire  _GEN_157; // @[mmu_conv.scala 109:45]
  wire  hit_12; // @[mmu_conv.scala 119:32]
  wire  _GEN_159; // @[mmu_conv.scala 126:35]
  wire  _GEN_160; // @[mmu_conv.scala 129:35]
  wire  _GEN_161; // @[mmu_conv.scala 130:35]
  wire  _T_427; // @[mmu_conv.scala 134:36]
  wire  _GEN_162; // @[mmu_conv.scala 134:61]
  wire  _GEN_163; // @[mmu_conv.scala 138:36]
  wire  _GEN_164; // @[mmu_conv.scala 133:21]
  wire  _GEN_165; // @[mmu_conv.scala 128:42]
  wire  protect_exception_12; // @[mmu_conv.scala 125:18]
  wire  _GEN_167; // @[mmu_conv.scala 145:32]
  wire  _T_436; // @[mmu_conv.scala 148:36]
  wire  update_exception_12; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_437; // @[Cat.scala 29:58]
  wire [33:0] _GEN_310; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_438; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_440; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_311; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_444; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_445; // @[mmu_conv.scala 113:64]
  wire  _T_446; // @[mmu_conv.scala 113:48]
  wire  _GEN_169; // @[mmu_conv.scala 112:50]
  wire  _GEN_170; // @[mmu_conv.scala 109:45]
  wire  hit_13; // @[mmu_conv.scala 119:32]
  wire  _GEN_172; // @[mmu_conv.scala 126:35]
  wire  _GEN_173; // @[mmu_conv.scala 129:35]
  wire  _GEN_174; // @[mmu_conv.scala 130:35]
  wire  _T_461; // @[mmu_conv.scala 134:36]
  wire  _GEN_175; // @[mmu_conv.scala 134:61]
  wire  _GEN_176; // @[mmu_conv.scala 138:36]
  wire  _GEN_177; // @[mmu_conv.scala 133:21]
  wire  _GEN_178; // @[mmu_conv.scala 128:42]
  wire  protect_exception_13; // @[mmu_conv.scala 125:18]
  wire  _GEN_180; // @[mmu_conv.scala 145:32]
  wire  _T_470; // @[mmu_conv.scala 148:36]
  wire  update_exception_13; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_471; // @[Cat.scala 29:58]
  wire [33:0] _GEN_312; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_472; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_474; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_313; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_478; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_479; // @[mmu_conv.scala 113:64]
  wire  _T_480; // @[mmu_conv.scala 113:48]
  wire  _GEN_182; // @[mmu_conv.scala 112:50]
  wire  _GEN_183; // @[mmu_conv.scala 109:45]
  wire  hit_14; // @[mmu_conv.scala 119:32]
  wire  _GEN_185; // @[mmu_conv.scala 126:35]
  wire  _GEN_186; // @[mmu_conv.scala 129:35]
  wire  _GEN_187; // @[mmu_conv.scala 130:35]
  wire  _T_495; // @[mmu_conv.scala 134:36]
  wire  _GEN_188; // @[mmu_conv.scala 134:61]
  wire  _GEN_189; // @[mmu_conv.scala 138:36]
  wire  _GEN_190; // @[mmu_conv.scala 133:21]
  wire  _GEN_191; // @[mmu_conv.scala 128:42]
  wire  protect_exception_14; // @[mmu_conv.scala 125:18]
  wire  _GEN_193; // @[mmu_conv.scala 145:32]
  wire  _T_504; // @[mmu_conv.scala 148:36]
  wire  update_exception_14; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_505; // @[Cat.scala 29:58]
  wire [33:0] _GEN_314; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_506; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_508; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_315; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_512; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_513; // @[mmu_conv.scala 113:64]
  wire  _T_514; // @[mmu_conv.scala 113:48]
  wire  _GEN_195; // @[mmu_conv.scala 112:50]
  wire  _GEN_196; // @[mmu_conv.scala 109:45]
  wire  hit_15; // @[mmu_conv.scala 119:32]
  wire  _GEN_198; // @[mmu_conv.scala 126:35]
  wire  _GEN_199; // @[mmu_conv.scala 129:35]
  wire  _GEN_200; // @[mmu_conv.scala 130:35]
  wire  _T_529; // @[mmu_conv.scala 134:36]
  wire  _GEN_201; // @[mmu_conv.scala 134:61]
  wire  _GEN_202; // @[mmu_conv.scala 138:36]
  wire  _GEN_203; // @[mmu_conv.scala 133:21]
  wire  _GEN_204; // @[mmu_conv.scala 128:42]
  wire  protect_exception_15; // @[mmu_conv.scala 125:18]
  wire  _GEN_206; // @[mmu_conv.scala 145:32]
  wire  _T_538; // @[mmu_conv.scala 148:36]
  wire  update_exception_15; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_539; // @[Cat.scala 29:58]
  wire [33:0] _GEN_316; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_540; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_542; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_317; // @[mmu_conv.scala 152:62]
  wire [7:0] _T_550; // @[mmu_conv.scala 158:33]
  wire [15:0] _T_558; // @[mmu_conv.scala 158:33]
  wire  _T_559; // @[mmu_conv.scala 158:40]
  wire  tlb_miss_exception; // @[mmu_conv.scala 158:28]
  wire [3:0] _GEN_208; // @[mmu_conv.scala 161:17]
  wire [3:0] _GEN_209; // @[mmu_conv.scala 162:17]
  wire [3:0] _GEN_210; // @[mmu_conv.scala 163:17]
  wire [3:0] _GEN_211; // @[mmu_conv.scala 164:17]
  wire [3:0] _GEN_212; // @[mmu_conv.scala 165:17]
  wire [3:0] _GEN_213; // @[mmu_conv.scala 166:17]
  wire [3:0] _GEN_214; // @[mmu_conv.scala 167:17]
  wire [3:0] _GEN_215; // @[mmu_conv.scala 168:17]
  wire [3:0] _GEN_216; // @[mmu_conv.scala 169:17]
  wire [3:0] _GEN_217; // @[mmu_conv.scala 170:17]
  wire [3:0] _GEN_218; // @[mmu_conv.scala 171:17]
  wire [3:0] _GEN_219; // @[mmu_conv.scala 172:17]
  wire [3:0] _GEN_220; // @[mmu_conv.scala 173:17]
  wire [3:0] _GEN_221; // @[mmu_conv.scala 174:17]
  wire [3:0] _GEN_222; // @[mmu_conv.scala 175:17]
  wire  _GEN_225; // @[mmu_conv.scala 178:39]
  wire  _GEN_226; // @[mmu_conv.scala 178:39]
  wire  _GEN_227; // @[mmu_conv.scala 178:39]
  wire  _GEN_228; // @[mmu_conv.scala 178:39]
  wire  _GEN_229; // @[mmu_conv.scala 178:39]
  wire  _GEN_230; // @[mmu_conv.scala 178:39]
  wire  _GEN_231; // @[mmu_conv.scala 178:39]
  wire  _GEN_232; // @[mmu_conv.scala 178:39]
  wire  _GEN_233; // @[mmu_conv.scala 178:39]
  wire  _GEN_234; // @[mmu_conv.scala 178:39]
  wire  _GEN_235; // @[mmu_conv.scala 178:39]
  wire  _GEN_236; // @[mmu_conv.scala 178:39]
  wire  _GEN_237; // @[mmu_conv.scala 178:39]
  wire  _GEN_238; // @[mmu_conv.scala 178:39]
  wire  _GEN_239; // @[mmu_conv.scala 178:39]
  wire  _T_562; // @[mmu_conv.scala 178:39]
  wire  _GEN_241; // @[mmu_conv.scala 178:75]
  wire  _GEN_242; // @[mmu_conv.scala 178:75]
  wire  _GEN_243; // @[mmu_conv.scala 178:75]
  wire  _GEN_244; // @[mmu_conv.scala 178:75]
  wire  _GEN_245; // @[mmu_conv.scala 178:75]
  wire  _GEN_246; // @[mmu_conv.scala 178:75]
  wire  _GEN_247; // @[mmu_conv.scala 178:75]
  wire  _GEN_248; // @[mmu_conv.scala 178:75]
  wire  _GEN_249; // @[mmu_conv.scala 178:75]
  wire  _GEN_250; // @[mmu_conv.scala 178:75]
  wire  _GEN_251; // @[mmu_conv.scala 178:75]
  wire  _GEN_252; // @[mmu_conv.scala 178:75]
  wire  _GEN_253; // @[mmu_conv.scala 178:75]
  wire  _GEN_254; // @[mmu_conv.scala 178:75]
  wire  _GEN_255; // @[mmu_conv.scala 178:75]
  wire  tlb_exception; // @[mmu_conv.scala 178:75]
  wire  _T_566; // @[mmu_conv.scala 191:23]
  wire  _T_568; // @[mmu_conv.scala 191:35]
  wire [33:0] _GEN_257; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_258; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_259; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_260; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_261; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_262; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_263; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_264; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_265; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_266; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_267; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_268; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_269; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_270; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_271; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_272; // @[mmu_conv.scala 200:36]
  wire  _GEN_273; // @[mmu_conv.scala 204:36]
  wire [33:0] _GEN_274; // @[mmu_conv.scala 198:48]
  wire  _GEN_275; // @[mmu_conv.scala 198:48]
  wire  _GEN_276; // @[mmu_conv.scala 198:48]
  wire [33:0] _GEN_277; // @[mmu_conv.scala 191:73]
  wire  _GEN_278; // @[mmu_conv.scala 191:73]
  wire  _GEN_279; // @[mmu_conv.scala 191:73]
  wire [33:0] _GEN_280; // @[mmu_conv.scala 186:40]
  wire  _GEN_281; // @[mmu_conv.scala 186:40]
  wire  _GEN_282; // @[mmu_conv.scala 186:40]
  assign _T = io_vm_i == 5'h0; // @[mmu_conv.scala 109:18]
  assign _T_1 = io_vm_i == 5'h8; // @[mmu_conv.scala 112:24]
  assign _T_2 = io_vir_addr_i & tlb_mask_0; // @[mmu_conv.scala 113:33]
  assign _T_3 = tlb_vpn_0 & tlb_mask_0; // @[mmu_conv.scala 113:64]
  assign _T_4 = _T_2 == _T_3; // @[mmu_conv.scala 113:48]
  assign _GEN_0 = _T_1 & _T_4; // @[mmu_conv.scala 112:50]
  assign _GEN_1 = _T ? 1'h0 : _GEN_0; // @[mmu_conv.scala 109:45]
  assign hit_0 = tlb_pte_0[0] ? _GEN_1 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_3 = ~tlb_pte_0[3] | ~hit_0; // @[mmu_conv.scala 126:35]
  assign _GEN_4 = ~tlb_pte_0[2] | ~hit_0; // @[mmu_conv.scala 129:35]
  assign _GEN_5 = ~tlb_pte_0[1] | _GEN_4; // @[mmu_conv.scala 130:35]
  assign _T_19 = ~tlb_pte_0[1] & ~tlb_pte_0[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_6 = _T_19 | ~hit_0; // @[mmu_conv.scala 134:61]
  assign _GEN_7 = ~tlb_pte_0[1] | ~hit_0; // @[mmu_conv.scala 138:36]
  assign _GEN_8 = io_mxr_i ? _GEN_6 : _GEN_7; // @[mmu_conv.scala 133:21]
  assign _GEN_9 = io_we_i ? _GEN_5 : _GEN_8; // @[mmu_conv.scala 128:42]
  assign protect_exception_0 = io_ex_i ? _GEN_3 : _GEN_9; // @[mmu_conv.scala 125:18]
  assign _GEN_11 = ~tlb_pte_0[6] | ~hit_0; // @[mmu_conv.scala 145:32]
  assign _T_28 = io_we_i & ~tlb_pte_0[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_0 = _T_28 | _GEN_11; // @[mmu_conv.scala 148:61]
  assign _T_29 = {tlb_pte_0,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_286 = {{2'd0}, tlb_mask_0}; // @[mmu_conv.scala 152:47]
  assign _T_30 = _T_29 & _GEN_286; // @[mmu_conv.scala 152:47]
  assign _T_32 = io_vir_addr_i & ~tlb_mask_0; // @[mmu_conv.scala 152:79]
  assign _GEN_287 = {{2'd0}, _T_32}; // @[mmu_conv.scala 152:62]
  assign _T_36 = io_vir_addr_i & tlb_mask_1; // @[mmu_conv.scala 113:33]
  assign _T_37 = tlb_vpn_1 & tlb_mask_1; // @[mmu_conv.scala 113:64]
  assign _T_38 = _T_36 == _T_37; // @[mmu_conv.scala 113:48]
  assign _GEN_13 = _T_1 & _T_38; // @[mmu_conv.scala 112:50]
  assign _GEN_14 = _T ? 1'h0 : _GEN_13; // @[mmu_conv.scala 109:45]
  assign hit_1 = tlb_pte_1[0] ? _GEN_14 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_16 = ~tlb_pte_1[3] | ~hit_1; // @[mmu_conv.scala 126:35]
  assign _GEN_17 = ~tlb_pte_1[2] | ~hit_1; // @[mmu_conv.scala 129:35]
  assign _GEN_18 = ~tlb_pte_1[1] | _GEN_17; // @[mmu_conv.scala 130:35]
  assign _T_53 = ~tlb_pte_1[1] & ~tlb_pte_1[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_19 = _T_53 | ~hit_1; // @[mmu_conv.scala 134:61]
  assign _GEN_20 = ~tlb_pte_1[1] | ~hit_1; // @[mmu_conv.scala 138:36]
  assign _GEN_21 = io_mxr_i ? _GEN_19 : _GEN_20; // @[mmu_conv.scala 133:21]
  assign _GEN_22 = io_we_i ? _GEN_18 : _GEN_21; // @[mmu_conv.scala 128:42]
  assign protect_exception_1 = io_ex_i ? _GEN_16 : _GEN_22; // @[mmu_conv.scala 125:18]
  assign _GEN_24 = ~tlb_pte_1[6] | ~hit_1; // @[mmu_conv.scala 145:32]
  assign _T_62 = io_we_i & ~tlb_pte_1[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_1 = _T_62 | _GEN_24; // @[mmu_conv.scala 148:61]
  assign _T_63 = {tlb_pte_1,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_288 = {{2'd0}, tlb_mask_1}; // @[mmu_conv.scala 152:47]
  assign _T_64 = _T_63 & _GEN_288; // @[mmu_conv.scala 152:47]
  assign _T_66 = io_vir_addr_i & ~tlb_mask_1; // @[mmu_conv.scala 152:79]
  assign _GEN_289 = {{2'd0}, _T_66}; // @[mmu_conv.scala 152:62]
  assign _T_70 = io_vir_addr_i & tlb_mask_2; // @[mmu_conv.scala 113:33]
  assign _T_71 = tlb_vpn_2 & tlb_mask_2; // @[mmu_conv.scala 113:64]
  assign _T_72 = _T_70 == _T_71; // @[mmu_conv.scala 113:48]
  assign _GEN_26 = _T_1 & _T_72; // @[mmu_conv.scala 112:50]
  assign _GEN_27 = _T ? 1'h0 : _GEN_26; // @[mmu_conv.scala 109:45]
  assign hit_2 = tlb_pte_2[0] ? _GEN_27 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_29 = ~tlb_pte_2[3] | ~hit_2; // @[mmu_conv.scala 126:35]
  assign _GEN_30 = ~tlb_pte_2[2] | ~hit_2; // @[mmu_conv.scala 129:35]
  assign _GEN_31 = ~tlb_pte_2[1] | _GEN_30; // @[mmu_conv.scala 130:35]
  assign _T_87 = ~tlb_pte_2[1] & ~tlb_pte_2[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_32 = _T_87 | ~hit_2; // @[mmu_conv.scala 134:61]
  assign _GEN_33 = ~tlb_pte_2[1] | ~hit_2; // @[mmu_conv.scala 138:36]
  assign _GEN_34 = io_mxr_i ? _GEN_32 : _GEN_33; // @[mmu_conv.scala 133:21]
  assign _GEN_35 = io_we_i ? _GEN_31 : _GEN_34; // @[mmu_conv.scala 128:42]
  assign protect_exception_2 = io_ex_i ? _GEN_29 : _GEN_35; // @[mmu_conv.scala 125:18]
  assign _GEN_37 = ~tlb_pte_2[6] | ~hit_2; // @[mmu_conv.scala 145:32]
  assign _T_96 = io_we_i & ~tlb_pte_2[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_2 = _T_96 | _GEN_37; // @[mmu_conv.scala 148:61]
  assign _T_97 = {tlb_pte_2,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_290 = {{2'd0}, tlb_mask_2}; // @[mmu_conv.scala 152:47]
  assign _T_98 = _T_97 & _GEN_290; // @[mmu_conv.scala 152:47]
  assign _T_100 = io_vir_addr_i & ~tlb_mask_2; // @[mmu_conv.scala 152:79]
  assign _GEN_291 = {{2'd0}, _T_100}; // @[mmu_conv.scala 152:62]
  assign _T_104 = io_vir_addr_i & tlb_mask_3; // @[mmu_conv.scala 113:33]
  assign _T_105 = tlb_vpn_3 & tlb_mask_3; // @[mmu_conv.scala 113:64]
  assign _T_106 = _T_104 == _T_105; // @[mmu_conv.scala 113:48]
  assign _GEN_39 = _T_1 & _T_106; // @[mmu_conv.scala 112:50]
  assign _GEN_40 = _T ? 1'h0 : _GEN_39; // @[mmu_conv.scala 109:45]
  assign hit_3 = tlb_pte_3[0] ? _GEN_40 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_42 = ~tlb_pte_3[3] | ~hit_3; // @[mmu_conv.scala 126:35]
  assign _GEN_43 = ~tlb_pte_3[2] | ~hit_3; // @[mmu_conv.scala 129:35]
  assign _GEN_44 = ~tlb_pte_3[1] | _GEN_43; // @[mmu_conv.scala 130:35]
  assign _T_121 = ~tlb_pte_3[1] & ~tlb_pte_3[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_45 = _T_121 | ~hit_3; // @[mmu_conv.scala 134:61]
  assign _GEN_46 = ~tlb_pte_3[1] | ~hit_3; // @[mmu_conv.scala 138:36]
  assign _GEN_47 = io_mxr_i ? _GEN_45 : _GEN_46; // @[mmu_conv.scala 133:21]
  assign _GEN_48 = io_we_i ? _GEN_44 : _GEN_47; // @[mmu_conv.scala 128:42]
  assign protect_exception_3 = io_ex_i ? _GEN_42 : _GEN_48; // @[mmu_conv.scala 125:18]
  assign _GEN_50 = ~tlb_pte_3[6] | ~hit_3; // @[mmu_conv.scala 145:32]
  assign _T_130 = io_we_i & ~tlb_pte_3[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_3 = _T_130 | _GEN_50; // @[mmu_conv.scala 148:61]
  assign _T_131 = {tlb_pte_3,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_292 = {{2'd0}, tlb_mask_3}; // @[mmu_conv.scala 152:47]
  assign _T_132 = _T_131 & _GEN_292; // @[mmu_conv.scala 152:47]
  assign _T_134 = io_vir_addr_i & ~tlb_mask_3; // @[mmu_conv.scala 152:79]
  assign _GEN_293 = {{2'd0}, _T_134}; // @[mmu_conv.scala 152:62]
  assign _T_138 = io_vir_addr_i & tlb_mask_4; // @[mmu_conv.scala 113:33]
  assign _T_139 = tlb_vpn_4 & tlb_mask_4; // @[mmu_conv.scala 113:64]
  assign _T_140 = _T_138 == _T_139; // @[mmu_conv.scala 113:48]
  assign _GEN_52 = _T_1 & _T_140; // @[mmu_conv.scala 112:50]
  assign _GEN_53 = _T ? 1'h0 : _GEN_52; // @[mmu_conv.scala 109:45]
  assign hit_4 = tlb_pte_4[0] ? _GEN_53 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_55 = ~tlb_pte_4[3] | ~hit_4; // @[mmu_conv.scala 126:35]
  assign _GEN_56 = ~tlb_pte_4[2] | ~hit_4; // @[mmu_conv.scala 129:35]
  assign _GEN_57 = ~tlb_pte_4[1] | _GEN_56; // @[mmu_conv.scala 130:35]
  assign _T_155 = ~tlb_pte_4[1] & ~tlb_pte_4[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_58 = _T_155 | ~hit_4; // @[mmu_conv.scala 134:61]
  assign _GEN_59 = ~tlb_pte_4[1] | ~hit_4; // @[mmu_conv.scala 138:36]
  assign _GEN_60 = io_mxr_i ? _GEN_58 : _GEN_59; // @[mmu_conv.scala 133:21]
  assign _GEN_61 = io_we_i ? _GEN_57 : _GEN_60; // @[mmu_conv.scala 128:42]
  assign protect_exception_4 = io_ex_i ? _GEN_55 : _GEN_61; // @[mmu_conv.scala 125:18]
  assign _GEN_63 = ~tlb_pte_4[6] | ~hit_4; // @[mmu_conv.scala 145:32]
  assign _T_164 = io_we_i & ~tlb_pte_4[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_4 = _T_164 | _GEN_63; // @[mmu_conv.scala 148:61]
  assign _T_165 = {tlb_pte_4,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_294 = {{2'd0}, tlb_mask_4}; // @[mmu_conv.scala 152:47]
  assign _T_166 = _T_165 & _GEN_294; // @[mmu_conv.scala 152:47]
  assign _T_168 = io_vir_addr_i & ~tlb_mask_4; // @[mmu_conv.scala 152:79]
  assign _GEN_295 = {{2'd0}, _T_168}; // @[mmu_conv.scala 152:62]
  assign _T_172 = io_vir_addr_i & tlb_mask_5; // @[mmu_conv.scala 113:33]
  assign _T_173 = tlb_vpn_5 & tlb_mask_5; // @[mmu_conv.scala 113:64]
  assign _T_174 = _T_172 == _T_173; // @[mmu_conv.scala 113:48]
  assign _GEN_65 = _T_1 & _T_174; // @[mmu_conv.scala 112:50]
  assign _GEN_66 = _T ? 1'h0 : _GEN_65; // @[mmu_conv.scala 109:45]
  assign hit_5 = tlb_pte_5[0] ? _GEN_66 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_68 = ~tlb_pte_5[3] | ~hit_5; // @[mmu_conv.scala 126:35]
  assign _GEN_69 = ~tlb_pte_5[2] | ~hit_5; // @[mmu_conv.scala 129:35]
  assign _GEN_70 = ~tlb_pte_5[1] | _GEN_69; // @[mmu_conv.scala 130:35]
  assign _T_189 = ~tlb_pte_5[1] & ~tlb_pte_5[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_71 = _T_189 | ~hit_5; // @[mmu_conv.scala 134:61]
  assign _GEN_72 = ~tlb_pte_5[1] | ~hit_5; // @[mmu_conv.scala 138:36]
  assign _GEN_73 = io_mxr_i ? _GEN_71 : _GEN_72; // @[mmu_conv.scala 133:21]
  assign _GEN_74 = io_we_i ? _GEN_70 : _GEN_73; // @[mmu_conv.scala 128:42]
  assign protect_exception_5 = io_ex_i ? _GEN_68 : _GEN_74; // @[mmu_conv.scala 125:18]
  assign _GEN_76 = ~tlb_pte_5[6] | ~hit_5; // @[mmu_conv.scala 145:32]
  assign _T_198 = io_we_i & ~tlb_pte_5[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_5 = _T_198 | _GEN_76; // @[mmu_conv.scala 148:61]
  assign _T_199 = {tlb_pte_5,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_296 = {{2'd0}, tlb_mask_5}; // @[mmu_conv.scala 152:47]
  assign _T_200 = _T_199 & _GEN_296; // @[mmu_conv.scala 152:47]
  assign _T_202 = io_vir_addr_i & ~tlb_mask_5; // @[mmu_conv.scala 152:79]
  assign _GEN_297 = {{2'd0}, _T_202}; // @[mmu_conv.scala 152:62]
  assign _T_206 = io_vir_addr_i & tlb_mask_6; // @[mmu_conv.scala 113:33]
  assign _T_207 = tlb_vpn_6 & tlb_mask_6; // @[mmu_conv.scala 113:64]
  assign _T_208 = _T_206 == _T_207; // @[mmu_conv.scala 113:48]
  assign _GEN_78 = _T_1 & _T_208; // @[mmu_conv.scala 112:50]
  assign _GEN_79 = _T ? 1'h0 : _GEN_78; // @[mmu_conv.scala 109:45]
  assign hit_6 = tlb_pte_6[0] ? _GEN_79 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_81 = ~tlb_pte_6[3] | ~hit_6; // @[mmu_conv.scala 126:35]
  assign _GEN_82 = ~tlb_pte_6[2] | ~hit_6; // @[mmu_conv.scala 129:35]
  assign _GEN_83 = ~tlb_pte_6[1] | _GEN_82; // @[mmu_conv.scala 130:35]
  assign _T_223 = ~tlb_pte_6[1] & ~tlb_pte_6[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_84 = _T_223 | ~hit_6; // @[mmu_conv.scala 134:61]
  assign _GEN_85 = ~tlb_pte_6[1] | ~hit_6; // @[mmu_conv.scala 138:36]
  assign _GEN_86 = io_mxr_i ? _GEN_84 : _GEN_85; // @[mmu_conv.scala 133:21]
  assign _GEN_87 = io_we_i ? _GEN_83 : _GEN_86; // @[mmu_conv.scala 128:42]
  assign protect_exception_6 = io_ex_i ? _GEN_81 : _GEN_87; // @[mmu_conv.scala 125:18]
  assign _GEN_89 = ~tlb_pte_6[6] | ~hit_6; // @[mmu_conv.scala 145:32]
  assign _T_232 = io_we_i & ~tlb_pte_6[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_6 = _T_232 | _GEN_89; // @[mmu_conv.scala 148:61]
  assign _T_233 = {tlb_pte_6,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_298 = {{2'd0}, tlb_mask_6}; // @[mmu_conv.scala 152:47]
  assign _T_234 = _T_233 & _GEN_298; // @[mmu_conv.scala 152:47]
  assign _T_236 = io_vir_addr_i & ~tlb_mask_6; // @[mmu_conv.scala 152:79]
  assign _GEN_299 = {{2'd0}, _T_236}; // @[mmu_conv.scala 152:62]
  assign _T_240 = io_vir_addr_i & tlb_mask_7; // @[mmu_conv.scala 113:33]
  assign _T_241 = tlb_vpn_7 & tlb_mask_7; // @[mmu_conv.scala 113:64]
  assign _T_242 = _T_240 == _T_241; // @[mmu_conv.scala 113:48]
  assign _GEN_91 = _T_1 & _T_242; // @[mmu_conv.scala 112:50]
  assign _GEN_92 = _T ? 1'h0 : _GEN_91; // @[mmu_conv.scala 109:45]
  assign hit_7 = tlb_pte_7[0] ? _GEN_92 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_94 = ~tlb_pte_7[3] | ~hit_7; // @[mmu_conv.scala 126:35]
  assign _GEN_95 = ~tlb_pte_7[2] | ~hit_7; // @[mmu_conv.scala 129:35]
  assign _GEN_96 = ~tlb_pte_7[1] | _GEN_95; // @[mmu_conv.scala 130:35]
  assign _T_257 = ~tlb_pte_7[1] & ~tlb_pte_7[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_97 = _T_257 | ~hit_7; // @[mmu_conv.scala 134:61]
  assign _GEN_98 = ~tlb_pte_7[1] | ~hit_7; // @[mmu_conv.scala 138:36]
  assign _GEN_99 = io_mxr_i ? _GEN_97 : _GEN_98; // @[mmu_conv.scala 133:21]
  assign _GEN_100 = io_we_i ? _GEN_96 : _GEN_99; // @[mmu_conv.scala 128:42]
  assign protect_exception_7 = io_ex_i ? _GEN_94 : _GEN_100; // @[mmu_conv.scala 125:18]
  assign _GEN_102 = ~tlb_pte_7[6] | ~hit_7; // @[mmu_conv.scala 145:32]
  assign _T_266 = io_we_i & ~tlb_pte_7[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_7 = _T_266 | _GEN_102; // @[mmu_conv.scala 148:61]
  assign _T_267 = {tlb_pte_7,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_300 = {{2'd0}, tlb_mask_7}; // @[mmu_conv.scala 152:47]
  assign _T_268 = _T_267 & _GEN_300; // @[mmu_conv.scala 152:47]
  assign _T_270 = io_vir_addr_i & ~tlb_mask_7; // @[mmu_conv.scala 152:79]
  assign _GEN_301 = {{2'd0}, _T_270}; // @[mmu_conv.scala 152:62]
  assign _T_274 = io_vir_addr_i & tlb_mask_8; // @[mmu_conv.scala 113:33]
  assign _T_275 = tlb_vpn_8 & tlb_mask_8; // @[mmu_conv.scala 113:64]
  assign _T_276 = _T_274 == _T_275; // @[mmu_conv.scala 113:48]
  assign _GEN_104 = _T_1 & _T_276; // @[mmu_conv.scala 112:50]
  assign _GEN_105 = _T ? 1'h0 : _GEN_104; // @[mmu_conv.scala 109:45]
  assign hit_8 = tlb_pte_8[0] ? _GEN_105 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_107 = ~tlb_pte_8[3] | ~hit_8; // @[mmu_conv.scala 126:35]
  assign _GEN_108 = ~tlb_pte_8[2] | ~hit_8; // @[mmu_conv.scala 129:35]
  assign _GEN_109 = ~tlb_pte_8[1] | _GEN_108; // @[mmu_conv.scala 130:35]
  assign _T_291 = ~tlb_pte_8[1] & ~tlb_pte_8[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_110 = _T_291 | ~hit_8; // @[mmu_conv.scala 134:61]
  assign _GEN_111 = ~tlb_pte_8[1] | ~hit_8; // @[mmu_conv.scala 138:36]
  assign _GEN_112 = io_mxr_i ? _GEN_110 : _GEN_111; // @[mmu_conv.scala 133:21]
  assign _GEN_113 = io_we_i ? _GEN_109 : _GEN_112; // @[mmu_conv.scala 128:42]
  assign protect_exception_8 = io_ex_i ? _GEN_107 : _GEN_113; // @[mmu_conv.scala 125:18]
  assign _GEN_115 = ~tlb_pte_8[6] | ~hit_8; // @[mmu_conv.scala 145:32]
  assign _T_300 = io_we_i & ~tlb_pte_8[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_8 = _T_300 | _GEN_115; // @[mmu_conv.scala 148:61]
  assign _T_301 = {tlb_pte_8,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_302 = {{2'd0}, tlb_mask_8}; // @[mmu_conv.scala 152:47]
  assign _T_302 = _T_301 & _GEN_302; // @[mmu_conv.scala 152:47]
  assign _T_304 = io_vir_addr_i & ~tlb_mask_8; // @[mmu_conv.scala 152:79]
  assign _GEN_303 = {{2'd0}, _T_304}; // @[mmu_conv.scala 152:62]
  assign _T_308 = io_vir_addr_i & tlb_mask_9; // @[mmu_conv.scala 113:33]
  assign _T_309 = tlb_vpn_9 & tlb_mask_9; // @[mmu_conv.scala 113:64]
  assign _T_310 = _T_308 == _T_309; // @[mmu_conv.scala 113:48]
  assign _GEN_117 = _T_1 & _T_310; // @[mmu_conv.scala 112:50]
  assign _GEN_118 = _T ? 1'h0 : _GEN_117; // @[mmu_conv.scala 109:45]
  assign hit_9 = tlb_pte_9[0] ? _GEN_118 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_120 = ~tlb_pte_9[3] | ~hit_9; // @[mmu_conv.scala 126:35]
  assign _GEN_121 = ~tlb_pte_9[2] | ~hit_9; // @[mmu_conv.scala 129:35]
  assign _GEN_122 = ~tlb_pte_9[1] | _GEN_121; // @[mmu_conv.scala 130:35]
  assign _T_325 = ~tlb_pte_9[1] & ~tlb_pte_9[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_123 = _T_325 | ~hit_9; // @[mmu_conv.scala 134:61]
  assign _GEN_124 = ~tlb_pte_9[1] | ~hit_9; // @[mmu_conv.scala 138:36]
  assign _GEN_125 = io_mxr_i ? _GEN_123 : _GEN_124; // @[mmu_conv.scala 133:21]
  assign _GEN_126 = io_we_i ? _GEN_122 : _GEN_125; // @[mmu_conv.scala 128:42]
  assign protect_exception_9 = io_ex_i ? _GEN_120 : _GEN_126; // @[mmu_conv.scala 125:18]
  assign _GEN_128 = ~tlb_pte_9[6] | ~hit_9; // @[mmu_conv.scala 145:32]
  assign _T_334 = io_we_i & ~tlb_pte_9[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_9 = _T_334 | _GEN_128; // @[mmu_conv.scala 148:61]
  assign _T_335 = {tlb_pte_9,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_304 = {{2'd0}, tlb_mask_9}; // @[mmu_conv.scala 152:47]
  assign _T_336 = _T_335 & _GEN_304; // @[mmu_conv.scala 152:47]
  assign _T_338 = io_vir_addr_i & ~tlb_mask_9; // @[mmu_conv.scala 152:79]
  assign _GEN_305 = {{2'd0}, _T_338}; // @[mmu_conv.scala 152:62]
  assign _T_342 = io_vir_addr_i & tlb_mask_10; // @[mmu_conv.scala 113:33]
  assign _T_343 = tlb_vpn_10 & tlb_mask_10; // @[mmu_conv.scala 113:64]
  assign _T_344 = _T_342 == _T_343; // @[mmu_conv.scala 113:48]
  assign _GEN_130 = _T_1 & _T_344; // @[mmu_conv.scala 112:50]
  assign _GEN_131 = _T ? 1'h0 : _GEN_130; // @[mmu_conv.scala 109:45]
  assign hit_10 = tlb_pte_10[0] ? _GEN_131 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_133 = ~tlb_pte_10[3] | ~hit_10; // @[mmu_conv.scala 126:35]
  assign _GEN_134 = ~tlb_pte_10[2] | ~hit_10; // @[mmu_conv.scala 129:35]
  assign _GEN_135 = ~tlb_pte_10[1] | _GEN_134; // @[mmu_conv.scala 130:35]
  assign _T_359 = ~tlb_pte_10[1] & ~tlb_pte_10[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_136 = _T_359 | ~hit_10; // @[mmu_conv.scala 134:61]
  assign _GEN_137 = ~tlb_pte_10[1] | ~hit_10; // @[mmu_conv.scala 138:36]
  assign _GEN_138 = io_mxr_i ? _GEN_136 : _GEN_137; // @[mmu_conv.scala 133:21]
  assign _GEN_139 = io_we_i ? _GEN_135 : _GEN_138; // @[mmu_conv.scala 128:42]
  assign protect_exception_10 = io_ex_i ? _GEN_133 : _GEN_139; // @[mmu_conv.scala 125:18]
  assign _GEN_141 = ~tlb_pte_10[6] | ~hit_10; // @[mmu_conv.scala 145:32]
  assign _T_368 = io_we_i & ~tlb_pte_10[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_10 = _T_368 | _GEN_141; // @[mmu_conv.scala 148:61]
  assign _T_369 = {tlb_pte_10,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_306 = {{2'd0}, tlb_mask_10}; // @[mmu_conv.scala 152:47]
  assign _T_370 = _T_369 & _GEN_306; // @[mmu_conv.scala 152:47]
  assign _T_372 = io_vir_addr_i & ~tlb_mask_10; // @[mmu_conv.scala 152:79]
  assign _GEN_307 = {{2'd0}, _T_372}; // @[mmu_conv.scala 152:62]
  assign _T_376 = io_vir_addr_i & tlb_mask_11; // @[mmu_conv.scala 113:33]
  assign _T_377 = tlb_vpn_11 & tlb_mask_11; // @[mmu_conv.scala 113:64]
  assign _T_378 = _T_376 == _T_377; // @[mmu_conv.scala 113:48]
  assign _GEN_143 = _T_1 & _T_378; // @[mmu_conv.scala 112:50]
  assign _GEN_144 = _T ? 1'h0 : _GEN_143; // @[mmu_conv.scala 109:45]
  assign hit_11 = tlb_pte_11[0] ? _GEN_144 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_146 = ~tlb_pte_11[3] | ~hit_11; // @[mmu_conv.scala 126:35]
  assign _GEN_147 = ~tlb_pte_11[2] | ~hit_11; // @[mmu_conv.scala 129:35]
  assign _GEN_148 = ~tlb_pte_11[1] | _GEN_147; // @[mmu_conv.scala 130:35]
  assign _T_393 = ~tlb_pte_11[1] & ~tlb_pte_11[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_149 = _T_393 | ~hit_11; // @[mmu_conv.scala 134:61]
  assign _GEN_150 = ~tlb_pte_11[1] | ~hit_11; // @[mmu_conv.scala 138:36]
  assign _GEN_151 = io_mxr_i ? _GEN_149 : _GEN_150; // @[mmu_conv.scala 133:21]
  assign _GEN_152 = io_we_i ? _GEN_148 : _GEN_151; // @[mmu_conv.scala 128:42]
  assign protect_exception_11 = io_ex_i ? _GEN_146 : _GEN_152; // @[mmu_conv.scala 125:18]
  assign _GEN_154 = ~tlb_pte_11[6] | ~hit_11; // @[mmu_conv.scala 145:32]
  assign _T_402 = io_we_i & ~tlb_pte_11[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_11 = _T_402 | _GEN_154; // @[mmu_conv.scala 148:61]
  assign _T_403 = {tlb_pte_11,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_308 = {{2'd0}, tlb_mask_11}; // @[mmu_conv.scala 152:47]
  assign _T_404 = _T_403 & _GEN_308; // @[mmu_conv.scala 152:47]
  assign _T_406 = io_vir_addr_i & ~tlb_mask_11; // @[mmu_conv.scala 152:79]
  assign _GEN_309 = {{2'd0}, _T_406}; // @[mmu_conv.scala 152:62]
  assign _T_410 = io_vir_addr_i & tlb_mask_12; // @[mmu_conv.scala 113:33]
  assign _T_411 = tlb_vpn_12 & tlb_mask_12; // @[mmu_conv.scala 113:64]
  assign _T_412 = _T_410 == _T_411; // @[mmu_conv.scala 113:48]
  assign _GEN_156 = _T_1 & _T_412; // @[mmu_conv.scala 112:50]
  assign _GEN_157 = _T ? 1'h0 : _GEN_156; // @[mmu_conv.scala 109:45]
  assign hit_12 = tlb_pte_12[0] ? _GEN_157 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_159 = ~tlb_pte_12[3] | ~hit_12; // @[mmu_conv.scala 126:35]
  assign _GEN_160 = ~tlb_pte_12[2] | ~hit_12; // @[mmu_conv.scala 129:35]
  assign _GEN_161 = ~tlb_pte_12[1] | _GEN_160; // @[mmu_conv.scala 130:35]
  assign _T_427 = ~tlb_pte_12[1] & ~tlb_pte_12[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_162 = _T_427 | ~hit_12; // @[mmu_conv.scala 134:61]
  assign _GEN_163 = ~tlb_pte_12[1] | ~hit_12; // @[mmu_conv.scala 138:36]
  assign _GEN_164 = io_mxr_i ? _GEN_162 : _GEN_163; // @[mmu_conv.scala 133:21]
  assign _GEN_165 = io_we_i ? _GEN_161 : _GEN_164; // @[mmu_conv.scala 128:42]
  assign protect_exception_12 = io_ex_i ? _GEN_159 : _GEN_165; // @[mmu_conv.scala 125:18]
  assign _GEN_167 = ~tlb_pte_12[6] | ~hit_12; // @[mmu_conv.scala 145:32]
  assign _T_436 = io_we_i & ~tlb_pte_12[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_12 = _T_436 | _GEN_167; // @[mmu_conv.scala 148:61]
  assign _T_437 = {tlb_pte_12,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_310 = {{2'd0}, tlb_mask_12}; // @[mmu_conv.scala 152:47]
  assign _T_438 = _T_437 & _GEN_310; // @[mmu_conv.scala 152:47]
  assign _T_440 = io_vir_addr_i & ~tlb_mask_12; // @[mmu_conv.scala 152:79]
  assign _GEN_311 = {{2'd0}, _T_440}; // @[mmu_conv.scala 152:62]
  assign _T_444 = io_vir_addr_i & tlb_mask_13; // @[mmu_conv.scala 113:33]
  assign _T_445 = tlb_vpn_13 & tlb_mask_13; // @[mmu_conv.scala 113:64]
  assign _T_446 = _T_444 == _T_445; // @[mmu_conv.scala 113:48]
  assign _GEN_169 = _T_1 & _T_446; // @[mmu_conv.scala 112:50]
  assign _GEN_170 = _T ? 1'h0 : _GEN_169; // @[mmu_conv.scala 109:45]
  assign hit_13 = tlb_pte_13[0] ? _GEN_170 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_172 = ~tlb_pte_13[3] | ~hit_13; // @[mmu_conv.scala 126:35]
  assign _GEN_173 = ~tlb_pte_13[2] | ~hit_13; // @[mmu_conv.scala 129:35]
  assign _GEN_174 = ~tlb_pte_13[1] | _GEN_173; // @[mmu_conv.scala 130:35]
  assign _T_461 = ~tlb_pte_13[1] & ~tlb_pte_13[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_175 = _T_461 | ~hit_13; // @[mmu_conv.scala 134:61]
  assign _GEN_176 = ~tlb_pte_13[1] | ~hit_13; // @[mmu_conv.scala 138:36]
  assign _GEN_177 = io_mxr_i ? _GEN_175 : _GEN_176; // @[mmu_conv.scala 133:21]
  assign _GEN_178 = io_we_i ? _GEN_174 : _GEN_177; // @[mmu_conv.scala 128:42]
  assign protect_exception_13 = io_ex_i ? _GEN_172 : _GEN_178; // @[mmu_conv.scala 125:18]
  assign _GEN_180 = ~tlb_pte_13[6] | ~hit_13; // @[mmu_conv.scala 145:32]
  assign _T_470 = io_we_i & ~tlb_pte_13[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_13 = _T_470 | _GEN_180; // @[mmu_conv.scala 148:61]
  assign _T_471 = {tlb_pte_13,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_312 = {{2'd0}, tlb_mask_13}; // @[mmu_conv.scala 152:47]
  assign _T_472 = _T_471 & _GEN_312; // @[mmu_conv.scala 152:47]
  assign _T_474 = io_vir_addr_i & ~tlb_mask_13; // @[mmu_conv.scala 152:79]
  assign _GEN_313 = {{2'd0}, _T_474}; // @[mmu_conv.scala 152:62]
  assign _T_478 = io_vir_addr_i & tlb_mask_14; // @[mmu_conv.scala 113:33]
  assign _T_479 = tlb_vpn_14 & tlb_mask_14; // @[mmu_conv.scala 113:64]
  assign _T_480 = _T_478 == _T_479; // @[mmu_conv.scala 113:48]
  assign _GEN_182 = _T_1 & _T_480; // @[mmu_conv.scala 112:50]
  assign _GEN_183 = _T ? 1'h0 : _GEN_182; // @[mmu_conv.scala 109:45]
  assign hit_14 = tlb_pte_14[0] ? _GEN_183 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_185 = ~tlb_pte_14[3] | ~hit_14; // @[mmu_conv.scala 126:35]
  assign _GEN_186 = ~tlb_pte_14[2] | ~hit_14; // @[mmu_conv.scala 129:35]
  assign _GEN_187 = ~tlb_pte_14[1] | _GEN_186; // @[mmu_conv.scala 130:35]
  assign _T_495 = ~tlb_pte_14[1] & ~tlb_pte_14[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_188 = _T_495 | ~hit_14; // @[mmu_conv.scala 134:61]
  assign _GEN_189 = ~tlb_pte_14[1] | ~hit_14; // @[mmu_conv.scala 138:36]
  assign _GEN_190 = io_mxr_i ? _GEN_188 : _GEN_189; // @[mmu_conv.scala 133:21]
  assign _GEN_191 = io_we_i ? _GEN_187 : _GEN_190; // @[mmu_conv.scala 128:42]
  assign protect_exception_14 = io_ex_i ? _GEN_185 : _GEN_191; // @[mmu_conv.scala 125:18]
  assign _GEN_193 = ~tlb_pte_14[6] | ~hit_14; // @[mmu_conv.scala 145:32]
  assign _T_504 = io_we_i & ~tlb_pte_14[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_14 = _T_504 | _GEN_193; // @[mmu_conv.scala 148:61]
  assign _T_505 = {tlb_pte_14,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_314 = {{2'd0}, tlb_mask_14}; // @[mmu_conv.scala 152:47]
  assign _T_506 = _T_505 & _GEN_314; // @[mmu_conv.scala 152:47]
  assign _T_508 = io_vir_addr_i & ~tlb_mask_14; // @[mmu_conv.scala 152:79]
  assign _GEN_315 = {{2'd0}, _T_508}; // @[mmu_conv.scala 152:62]
  assign _T_512 = io_vir_addr_i & tlb_mask_15; // @[mmu_conv.scala 113:33]
  assign _T_513 = tlb_vpn_15 & tlb_mask_15; // @[mmu_conv.scala 113:64]
  assign _T_514 = _T_512 == _T_513; // @[mmu_conv.scala 113:48]
  assign _GEN_195 = _T_1 & _T_514; // @[mmu_conv.scala 112:50]
  assign _GEN_196 = _T ? 1'h0 : _GEN_195; // @[mmu_conv.scala 109:45]
  assign hit_15 = tlb_pte_15[0] ? _GEN_196 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_198 = ~tlb_pte_15[3] | ~hit_15; // @[mmu_conv.scala 126:35]
  assign _GEN_199 = ~tlb_pte_15[2] | ~hit_15; // @[mmu_conv.scala 129:35]
  assign _GEN_200 = ~tlb_pte_15[1] | _GEN_199; // @[mmu_conv.scala 130:35]
  assign _T_529 = ~tlb_pte_15[1] & ~tlb_pte_15[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_201 = _T_529 | ~hit_15; // @[mmu_conv.scala 134:61]
  assign _GEN_202 = ~tlb_pte_15[1] | ~hit_15; // @[mmu_conv.scala 138:36]
  assign _GEN_203 = io_mxr_i ? _GEN_201 : _GEN_202; // @[mmu_conv.scala 133:21]
  assign _GEN_204 = io_we_i ? _GEN_200 : _GEN_203; // @[mmu_conv.scala 128:42]
  assign protect_exception_15 = io_ex_i ? _GEN_198 : _GEN_204; // @[mmu_conv.scala 125:18]
  assign _GEN_206 = ~tlb_pte_15[6] | ~hit_15; // @[mmu_conv.scala 145:32]
  assign _T_538 = io_we_i & ~tlb_pte_15[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_15 = _T_538 | _GEN_206; // @[mmu_conv.scala 148:61]
  assign _T_539 = {tlb_pte_15,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_316 = {{2'd0}, tlb_mask_15}; // @[mmu_conv.scala 152:47]
  assign _T_540 = _T_539 & _GEN_316; // @[mmu_conv.scala 152:47]
  assign _T_542 = io_vir_addr_i & ~tlb_mask_15; // @[mmu_conv.scala 152:79]
  assign _GEN_317 = {{2'd0}, _T_542}; // @[mmu_conv.scala 152:62]
  assign _T_550 = {hit_7,hit_6,hit_5,hit_4,hit_3,hit_2,hit_1,hit_0}; // @[mmu_conv.scala 158:33]
  assign _T_558 = {hit_15,hit_14,hit_13,hit_12,hit_11,hit_10,hit_9,hit_8,_T_550}; // @[mmu_conv.scala 158:33]
  assign _T_559 = _T_558 != 16'h0; // @[mmu_conv.scala 158:40]
  assign tlb_miss_exception = _T_559 ? 1'h0 : 1'h1; // @[mmu_conv.scala 158:28]
  assign _GEN_208 = hit_15 ? 4'hf : 4'h0; // @[mmu_conv.scala 161:17]
  assign _GEN_209 = hit_14 ? 4'he : _GEN_208; // @[mmu_conv.scala 162:17]
  assign _GEN_210 = hit_13 ? 4'hd : _GEN_209; // @[mmu_conv.scala 163:17]
  assign _GEN_211 = hit_12 ? 4'hc : _GEN_210; // @[mmu_conv.scala 164:17]
  assign _GEN_212 = hit_11 ? 4'hb : _GEN_211; // @[mmu_conv.scala 165:17]
  assign _GEN_213 = hit_10 ? 4'ha : _GEN_212; // @[mmu_conv.scala 166:17]
  assign _GEN_214 = hit_9 ? 4'h9 : _GEN_213; // @[mmu_conv.scala 167:17]
  assign _GEN_215 = hit_8 ? 4'h8 : _GEN_214; // @[mmu_conv.scala 168:17]
  assign _GEN_216 = hit_7 ? 4'h7 : _GEN_215; // @[mmu_conv.scala 169:17]
  assign _GEN_217 = hit_6 ? 4'h6 : _GEN_216; // @[mmu_conv.scala 170:17]
  assign _GEN_218 = hit_5 ? 4'h5 : _GEN_217; // @[mmu_conv.scala 171:17]
  assign _GEN_219 = hit_4 ? 4'h4 : _GEN_218; // @[mmu_conv.scala 172:17]
  assign _GEN_220 = hit_3 ? 4'h3 : _GEN_219; // @[mmu_conv.scala 173:17]
  assign _GEN_221 = hit_2 ? 4'h2 : _GEN_220; // @[mmu_conv.scala 174:17]
  assign _GEN_222 = hit_1 ? 4'h1 : _GEN_221; // @[mmu_conv.scala 175:17]
  assign _GEN_225 = 4'h1 == io_hit_index_o ? protect_exception_1 : protect_exception_0; // @[mmu_conv.scala 178:39]
  assign _GEN_226 = 4'h2 == io_hit_index_o ? protect_exception_2 : _GEN_225; // @[mmu_conv.scala 178:39]
  assign _GEN_227 = 4'h3 == io_hit_index_o ? protect_exception_3 : _GEN_226; // @[mmu_conv.scala 178:39]
  assign _GEN_228 = 4'h4 == io_hit_index_o ? protect_exception_4 : _GEN_227; // @[mmu_conv.scala 178:39]
  assign _GEN_229 = 4'h5 == io_hit_index_o ? protect_exception_5 : _GEN_228; // @[mmu_conv.scala 178:39]
  assign _GEN_230 = 4'h6 == io_hit_index_o ? protect_exception_6 : _GEN_229; // @[mmu_conv.scala 178:39]
  assign _GEN_231 = 4'h7 == io_hit_index_o ? protect_exception_7 : _GEN_230; // @[mmu_conv.scala 178:39]
  assign _GEN_232 = 4'h8 == io_hit_index_o ? protect_exception_8 : _GEN_231; // @[mmu_conv.scala 178:39]
  assign _GEN_233 = 4'h9 == io_hit_index_o ? protect_exception_9 : _GEN_232; // @[mmu_conv.scala 178:39]
  assign _GEN_234 = 4'ha == io_hit_index_o ? protect_exception_10 : _GEN_233; // @[mmu_conv.scala 178:39]
  assign _GEN_235 = 4'hb == io_hit_index_o ? protect_exception_11 : _GEN_234; // @[mmu_conv.scala 178:39]
  assign _GEN_236 = 4'hc == io_hit_index_o ? protect_exception_12 : _GEN_235; // @[mmu_conv.scala 178:39]
  assign _GEN_237 = 4'hd == io_hit_index_o ? protect_exception_13 : _GEN_236; // @[mmu_conv.scala 178:39]
  assign _GEN_238 = 4'he == io_hit_index_o ? protect_exception_14 : _GEN_237; // @[mmu_conv.scala 178:39]
  assign _GEN_239 = 4'hf == io_hit_index_o ? protect_exception_15 : _GEN_238; // @[mmu_conv.scala 178:39]
  assign _T_562 = tlb_miss_exception | _GEN_239; // @[mmu_conv.scala 178:39]
  assign _GEN_241 = 4'h1 == io_hit_index_o ? update_exception_1 : update_exception_0; // @[mmu_conv.scala 178:75]
  assign _GEN_242 = 4'h2 == io_hit_index_o ? update_exception_2 : _GEN_241; // @[mmu_conv.scala 178:75]
  assign _GEN_243 = 4'h3 == io_hit_index_o ? update_exception_3 : _GEN_242; // @[mmu_conv.scala 178:75]
  assign _GEN_244 = 4'h4 == io_hit_index_o ? update_exception_4 : _GEN_243; // @[mmu_conv.scala 178:75]
  assign _GEN_245 = 4'h5 == io_hit_index_o ? update_exception_5 : _GEN_244; // @[mmu_conv.scala 178:75]
  assign _GEN_246 = 4'h6 == io_hit_index_o ? update_exception_6 : _GEN_245; // @[mmu_conv.scala 178:75]
  assign _GEN_247 = 4'h7 == io_hit_index_o ? update_exception_7 : _GEN_246; // @[mmu_conv.scala 178:75]
  assign _GEN_248 = 4'h8 == io_hit_index_o ? update_exception_8 : _GEN_247; // @[mmu_conv.scala 178:75]
  assign _GEN_249 = 4'h9 == io_hit_index_o ? update_exception_9 : _GEN_248; // @[mmu_conv.scala 178:75]
  assign _GEN_250 = 4'ha == io_hit_index_o ? update_exception_10 : _GEN_249; // @[mmu_conv.scala 178:75]
  assign _GEN_251 = 4'hb == io_hit_index_o ? update_exception_11 : _GEN_250; // @[mmu_conv.scala 178:75]
  assign _GEN_252 = 4'hc == io_hit_index_o ? update_exception_12 : _GEN_251; // @[mmu_conv.scala 178:75]
  assign _GEN_253 = 4'hd == io_hit_index_o ? update_exception_13 : _GEN_252; // @[mmu_conv.scala 178:75]
  assign _GEN_254 = 4'he == io_hit_index_o ? update_exception_14 : _GEN_253; // @[mmu_conv.scala 178:75]
  assign _GEN_255 = 4'hf == io_hit_index_o ? update_exception_15 : _GEN_254; // @[mmu_conv.scala 178:75]
  assign tlb_exception = _T_562 | _GEN_255; // @[mmu_conv.scala 178:75]
  assign _T_566 = io_prv_i == 2'h3; // @[mmu_conv.scala 191:23]
  assign _T_568 = _T_566 | _T; // @[mmu_conv.scala 191:35]
  assign _GEN_257 = 4'h1 == io_hit_index_o ? phy_addr_1 : phy_addr_0; // @[mmu_conv.scala 201:21]
  assign _GEN_258 = 4'h2 == io_hit_index_o ? phy_addr_2 : _GEN_257; // @[mmu_conv.scala 201:21]
  assign _GEN_259 = 4'h3 == io_hit_index_o ? phy_addr_3 : _GEN_258; // @[mmu_conv.scala 201:21]
  assign _GEN_260 = 4'h4 == io_hit_index_o ? phy_addr_4 : _GEN_259; // @[mmu_conv.scala 201:21]
  assign _GEN_261 = 4'h5 == io_hit_index_o ? phy_addr_5 : _GEN_260; // @[mmu_conv.scala 201:21]
  assign _GEN_262 = 4'h6 == io_hit_index_o ? phy_addr_6 : _GEN_261; // @[mmu_conv.scala 201:21]
  assign _GEN_263 = 4'h7 == io_hit_index_o ? phy_addr_7 : _GEN_262; // @[mmu_conv.scala 201:21]
  assign _GEN_264 = 4'h8 == io_hit_index_o ? phy_addr_8 : _GEN_263; // @[mmu_conv.scala 201:21]
  assign _GEN_265 = 4'h9 == io_hit_index_o ? phy_addr_9 : _GEN_264; // @[mmu_conv.scala 201:21]
  assign _GEN_266 = 4'ha == io_hit_index_o ? phy_addr_10 : _GEN_265; // @[mmu_conv.scala 201:21]
  assign _GEN_267 = 4'hb == io_hit_index_o ? phy_addr_11 : _GEN_266; // @[mmu_conv.scala 201:21]
  assign _GEN_268 = 4'hc == io_hit_index_o ? phy_addr_12 : _GEN_267; // @[mmu_conv.scala 201:21]
  assign _GEN_269 = 4'hd == io_hit_index_o ? phy_addr_13 : _GEN_268; // @[mmu_conv.scala 201:21]
  assign _GEN_270 = 4'he == io_hit_index_o ? phy_addr_14 : _GEN_269; // @[mmu_conv.scala 201:21]
  assign _GEN_271 = 4'hf == io_hit_index_o ? phy_addr_15 : _GEN_270; // @[mmu_conv.scala 201:21]
  assign _GEN_272 = tlb_exception ? 34'h0 : _GEN_271; // @[mmu_conv.scala 200:36]
  assign _GEN_273 = tlb_miss_exception ? 1'h0 : _GEN_255; // @[mmu_conv.scala 204:36]
  assign _GEN_274 = _T_1 ? _GEN_272 : 34'h0; // @[mmu_conv.scala 198:48]
  assign _GEN_275 = _T_1 & tlb_exception; // @[mmu_conv.scala 198:48]
  assign _GEN_276 = _T_1 & _GEN_273; // @[mmu_conv.scala 198:48]
  assign _GEN_277 = _T_568 ? {{2'd0}, io_vir_addr_i} : _GEN_274; // @[mmu_conv.scala 191:73]
  assign _GEN_278 = _T_568 ? 1'h0 : _GEN_275; // @[mmu_conv.scala 191:73]
  assign _GEN_279 = _T_568 ? 1'h0 : _GEN_276; // @[mmu_conv.scala 191:73]
  assign _GEN_280 = io_ce_i ? _GEN_277 : 34'h0; // @[mmu_conv.scala 186:40]
  assign _GEN_281 = io_ce_i ? _GEN_278 : 1'h0; // @[mmu_conv.scala 186:40]
  assign _GEN_282 = io_ce_i ? _GEN_279 : 1'h0; // @[mmu_conv.scala 186:40]
  assign io_phy_addr_o = io_rst_n ? _GEN_280 : 34'h0; // @[mmu_conv.scala 182:19 mmu_conv.scala 187:19 mmu_conv.scala 192:19 mmu_conv.scala 193:19 mmu_conv.scala 199:19 mmu_conv.scala 201:21 mmu_conv.scala 211:19]
  assign io_tlb_exception_o = io_rst_n ? _GEN_281 : 1'h0; // @[mmu_conv.scala 183:24 mmu_conv.scala 188:24 mmu_conv.scala 195:24 mmu_conv.scala 203:24 mmu_conv.scala 212:24]
  assign io_tlb_update_o = io_rst_n ? _GEN_282 : 1'h0; // @[mmu_conv.scala 184:21 mmu_conv.scala 189:21 mmu_conv.scala 196:21 mmu_conv.scala 205:23 mmu_conv.scala 207:23 mmu_conv.scala 213:21]
  assign io_hit_index_o = hit_0 ? 4'h0 : _GEN_222; // @[mmu_conv.scala 160:18 mmu_conv.scala 161:33 mmu_conv.scala 162:33 mmu_conv.scala 163:33 mmu_conv.scala 164:33 mmu_conv.scala 165:33 mmu_conv.scala 166:33 mmu_conv.scala 167:33 mmu_conv.scala 168:33 mmu_conv.scala 169:33 mmu_conv.scala 170:33 mmu_conv.scala 171:33 mmu_conv.scala 172:33 mmu_conv.scala 173:33 mmu_conv.scala 174:33 mmu_conv.scala 175:33 mmu_conv.scala 176:33]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tlb_vpn_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tlb_vpn_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  tlb_vpn_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  tlb_vpn_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  tlb_vpn_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  tlb_vpn_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  tlb_vpn_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  tlb_vpn_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tlb_vpn_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  tlb_vpn_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  tlb_vpn_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  tlb_vpn_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  tlb_vpn_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  tlb_vpn_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  tlb_vpn_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  tlb_vpn_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  tlb_pte_0 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  tlb_pte_1 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  tlb_pte_2 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  tlb_pte_3 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  tlb_pte_4 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  tlb_pte_5 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  tlb_pte_6 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  tlb_pte_7 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  tlb_pte_8 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  tlb_pte_9 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  tlb_pte_10 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  tlb_pte_11 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  tlb_pte_12 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  tlb_pte_13 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  tlb_pte_14 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  tlb_pte_15 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  tlb_mask_0 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  tlb_mask_1 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  tlb_mask_2 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  tlb_mask_3 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  tlb_mask_4 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  tlb_mask_5 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  tlb_mask_6 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  tlb_mask_7 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  tlb_mask_8 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  tlb_mask_9 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  tlb_mask_10 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  tlb_mask_11 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  tlb_mask_12 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  tlb_mask_13 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  tlb_mask_14 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  tlb_mask_15 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  phy_addr_0 = _RAND_48[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  phy_addr_1 = _RAND_49[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {2{`RANDOM}};
  phy_addr_2 = _RAND_50[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {2{`RANDOM}};
  phy_addr_3 = _RAND_51[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {2{`RANDOM}};
  phy_addr_4 = _RAND_52[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {2{`RANDOM}};
  phy_addr_5 = _RAND_53[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {2{`RANDOM}};
  phy_addr_6 = _RAND_54[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  phy_addr_7 = _RAND_55[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {2{`RANDOM}};
  phy_addr_8 = _RAND_56[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  phy_addr_9 = _RAND_57[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  phy_addr_10 = _RAND_58[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {2{`RANDOM}};
  phy_addr_11 = _RAND_59[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {2{`RANDOM}};
  phy_addr_12 = _RAND_60[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {2{`RANDOM}};
  phy_addr_13 = _RAND_61[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {2{`RANDOM}};
  phy_addr_14 = _RAND_62[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {2{`RANDOM}};
  phy_addr_15 = _RAND_63[33:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(*) begin
    tlb_vpn_0 <= io_tlb0_vpn_i;
    tlb_vpn_1 <= io_tlb1_vpn_i;
    tlb_vpn_2 <= io_tlb2_vpn_i;
    tlb_vpn_3 <= io_tlb3_vpn_i;
    tlb_vpn_4 <= io_tlb4_vpn_i;
    tlb_vpn_5 <= io_tlb5_vpn_i;
    tlb_vpn_6 <= io_tlb6_vpn_i;
    tlb_vpn_7 <= io_tlb7_vpn_i;
    tlb_vpn_8 <= io_tlb8_vpn_i;
    tlb_vpn_9 <= io_tlb9_vpn_i;
    tlb_vpn_10 <= io_tlb10_vpn_i;
    tlb_vpn_11 <= io_tlb11_vpn_i;
    tlb_vpn_12 <= io_tlb12_vpn_i;
    tlb_vpn_13 <= io_tlb13_vpn_i;
    tlb_vpn_14 <= io_tlb14_vpn_i;
    tlb_vpn_15 <= io_tlb15_vpn_i;
    tlb_pte_0 <= io_tlb0_pte_i;
    tlb_pte_1 <= io_tlb1_pte_i;
    tlb_pte_2 <= io_tlb2_pte_i;
    tlb_pte_3 <= io_tlb3_pte_i;
    tlb_pte_4 <= io_tlb4_pte_i;
    tlb_pte_5 <= io_tlb5_pte_i;
    tlb_pte_6 <= io_tlb6_pte_i;
    tlb_pte_7 <= io_tlb7_pte_i;
    tlb_pte_8 <= io_tlb8_pte_i;
    tlb_pte_9 <= io_tlb9_pte_i;
    tlb_pte_10 <= io_tlb10_pte_i;
    tlb_pte_11 <= io_tlb11_pte_i;
    tlb_pte_12 <= io_tlb12_pte_i;
    tlb_pte_13 <= io_tlb13_pte_i;
    tlb_pte_14 <= io_tlb14_pte_i;
    tlb_pte_15 <= io_tlb15_pte_i;
    tlb_mask_0 <= io_tlb0_mask_i;
    tlb_mask_1 <= io_tlb1_mask_i;
    tlb_mask_2 <= io_tlb2_mask_i;
    tlb_mask_3 <= io_tlb3_mask_i;
    tlb_mask_4 <= io_tlb4_mask_i;
    tlb_mask_5 <= io_tlb5_mask_i;
    tlb_mask_6 <= io_tlb6_mask_i;
    tlb_mask_7 <= io_tlb7_mask_i;
    tlb_mask_8 <= io_tlb8_mask_i;
    tlb_mask_9 <= io_tlb9_mask_i;
    tlb_mask_10 <= io_tlb10_mask_i;
    tlb_mask_11 <= io_tlb11_mask_i;
    tlb_mask_12 <= io_tlb12_mask_i;
    tlb_mask_13 <= io_tlb13_mask_i;
    tlb_mask_14 <= io_tlb14_mask_i;
    tlb_mask_15 <= io_tlb15_mask_i;
    phy_addr_0 <= _T_30 | _GEN_287;
    phy_addr_1 <= _T_64 | _GEN_289;
    phy_addr_2 <= _T_98 | _GEN_291;
    phy_addr_3 <= _T_132 | _GEN_293;
    phy_addr_4 <= _T_166 | _GEN_295;
    phy_addr_5 <= _T_200 | _GEN_297;
    phy_addr_6 <= _T_234 | _GEN_299;
    phy_addr_7 <= _T_268 | _GEN_301;
    phy_addr_8 <= _T_302 | _GEN_303;
    phy_addr_9 <= _T_336 | _GEN_305;
    phy_addr_10 <= _T_370 | _GEN_307;
    phy_addr_11 <= _T_404 | _GEN_309;
    phy_addr_12 <= _T_438 | _GEN_311;
    phy_addr_13 <= _T_472 | _GEN_313;
    phy_addr_14 <= _T_506 | _GEN_315;
    phy_addr_15 <= _T_540 | _GEN_317;
  end
endmodule
