module mmu_conv(
  input         io_rst_n,
  input  [31:0] io_tlb0_vpn_i,
  input  [31:0] io_tlb0_mask_i,
  input  [31:0] io_tlb0_pte_i,
  input  [31:0] io_tlb1_vpn_i,
  input  [31:0] io_tlb1_mask_i,
  input  [31:0] io_tlb1_pte_i,
  input  [31:0] io_tlb2_vpn_i,
  input  [31:0] io_tlb2_mask_i,
  input  [31:0] io_tlb2_pte_i,
  input  [31:0] io_tlb3_vpn_i,
  input  [31:0] io_tlb3_mask_i,
  input  [31:0] io_tlb3_pte_i,
  input  [31:0] io_tlb4_vpn_i,
  input  [31:0] io_tlb4_mask_i,
  input  [31:0] io_tlb4_pte_i,
  input  [31:0] io_tlb5_vpn_i,
  input  [31:0] io_tlb5_mask_i,
  input  [31:0] io_tlb5_pte_i,
  input  [31:0] io_tlb6_vpn_i,
  input  [31:0] io_tlb6_mask_i,
  input  [31:0] io_tlb6_pte_i,
  input  [31:0] io_tlb7_vpn_i,
  input  [31:0] io_tlb7_mask_i,
  input  [31:0] io_tlb7_pte_i,
  input  [31:0] io_tlb8_vpn_i,
  input  [31:0] io_tlb8_mask_i,
  input  [31:0] io_tlb8_pte_i,
  input  [31:0] io_tlb9_vpn_i,
  input  [31:0] io_tlb9_mask_i,
  input  [31:0] io_tlb9_pte_i,
  input  [31:0] io_tlb10_vpn_i,
  input  [31:0] io_tlb10_mask_i,
  input  [31:0] io_tlb10_pte_i,
  input  [31:0] io_tlb11_vpn_i,
  input  [31:0] io_tlb11_mask_i,
  input  [31:0] io_tlb11_pte_i,
  input  [31:0] io_tlb12_vpn_i,
  input  [31:0] io_tlb12_mask_i,
  input  [31:0] io_tlb12_pte_i,
  input  [31:0] io_tlb13_vpn_i,
  input  [31:0] io_tlb13_mask_i,
  input  [31:0] io_tlb13_pte_i,
  input  [31:0] io_tlb14_vpn_i,
  input  [31:0] io_tlb14_mask_i,
  input  [31:0] io_tlb14_pte_i,
  input  [31:0] io_tlb15_vpn_i,
  input  [31:0] io_tlb15_mask_i,
  input  [31:0] io_tlb15_pte_i,
  input  [4:0]  io_vm_i,
  input  [1:0]  io_prv_i,
  input         io_mxr_i,
  input         io_ce_i,
  input         io_ex_i,
  input         io_we_i,
  input  [31:0] io_vir_addr_i,
  output [33:0] io_phy_addr_o,
  output        io_tlb_exception_o,
  output        io_tlb_update_o,
  output [3:0]  io_hit_index_o
);
  reg [31:0] tlb_vpn_0; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_0;
  reg [31:0] tlb_vpn_1; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_1;
  reg [31:0] tlb_vpn_2; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_2;
  reg [31:0] tlb_vpn_3; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_3;
  reg [31:0] tlb_vpn_4; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_4;
  reg [31:0] tlb_vpn_5; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_5;
  reg [31:0] tlb_vpn_6; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_6;
  reg [31:0] tlb_vpn_7; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_7;
  reg [31:0] tlb_vpn_8; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_8;
  reg [31:0] tlb_vpn_9; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_9;
  reg [31:0] tlb_vpn_10; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_10;
  reg [31:0] tlb_vpn_11; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_11;
  reg [31:0] tlb_vpn_12; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_12;
  reg [31:0] tlb_vpn_13; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_13;
  reg [31:0] tlb_vpn_14; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_14;
  reg [31:0] tlb_vpn_15; // @[mmu_conv.scala 47:21]
  reg [31:0] _RAND_15;
  reg [31:0] tlb_pte_0; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_16;
  reg [31:0] tlb_pte_1; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_17;
  reg [31:0] tlb_pte_2; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_18;
  reg [31:0] tlb_pte_3; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_19;
  reg [31:0] tlb_pte_4; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_20;
  reg [31:0] tlb_pte_5; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_21;
  reg [31:0] tlb_pte_6; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_22;
  reg [31:0] tlb_pte_7; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_23;
  reg [31:0] tlb_pte_8; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_24;
  reg [31:0] tlb_pte_9; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_25;
  reg [31:0] tlb_pte_10; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_26;
  reg [31:0] tlb_pte_11; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_27;
  reg [31:0] tlb_pte_12; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_28;
  reg [31:0] tlb_pte_13; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_29;
  reg [31:0] tlb_pte_14; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_30;
  reg [31:0] tlb_pte_15; // @[mmu_conv.scala 48:21]
  reg [31:0] _RAND_31;
  reg [31:0] tlb_mask_0; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_32;
  reg [31:0] tlb_mask_1; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_33;
  reg [31:0] tlb_mask_2; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_34;
  reg [31:0] tlb_mask_3; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_35;
  reg [31:0] tlb_mask_4; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_36;
  reg [31:0] tlb_mask_5; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_37;
  reg [31:0] tlb_mask_6; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_38;
  reg [31:0] tlb_mask_7; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_39;
  reg [31:0] tlb_mask_8; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_40;
  reg [31:0] tlb_mask_9; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_41;
  reg [31:0] tlb_mask_10; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_42;
  reg [31:0] tlb_mask_11; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_43;
  reg [31:0] tlb_mask_12; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_44;
  reg [31:0] tlb_mask_13; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_45;
  reg [31:0] tlb_mask_14; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_46;
  reg [31:0] tlb_mask_15; // @[mmu_conv.scala 49:21]
  reg [31:0] _RAND_47;
  reg [33:0] phy_addr_0; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_48;
  reg [33:0] phy_addr_1; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_49;
  reg [33:0] phy_addr_2; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_50;
  reg [33:0] phy_addr_3; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_51;
  reg [33:0] phy_addr_4; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_52;
  reg [33:0] phy_addr_5; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_53;
  reg [33:0] phy_addr_6; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_54;
  reg [33:0] phy_addr_7; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_55;
  reg [33:0] phy_addr_8; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_56;
  reg [33:0] phy_addr_9; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_57;
  reg [33:0] phy_addr_10; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_58;
  reg [33:0] phy_addr_11; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_59;
  reg [33:0] phy_addr_12; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_60;
  reg [33:0] phy_addr_13; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_61;
  reg [33:0] phy_addr_14; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_62;
  reg [33:0] phy_addr_15; // @[mmu_conv.scala 106:21]
  reg [63:0] _RAND_63;
  wire  _T; // @[mmu_conv.scala 109:18]
  wire  _T_1; // @[mmu_conv.scala 112:24]
  wire [31:0] _T_2; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_3; // @[mmu_conv.scala 113:64]
  wire  _T_4; // @[mmu_conv.scala 113:48]
  wire  _GEN_0; // @[mmu_conv.scala 112:50]
  wire  _GEN_1; // @[mmu_conv.scala 109:45]
  wire  hit_0; // @[mmu_conv.scala 119:32]
  wire  _GEN_3; // @[mmu_conv.scala 126:35]
  wire  _GEN_4; // @[mmu_conv.scala 129:35]
  wire  _GEN_5; // @[mmu_conv.scala 130:35]
  wire  _T_19; // @[mmu_conv.scala 134:36]
  wire  _GEN_6; // @[mmu_conv.scala 134:61]
  wire  _GEN_7; // @[mmu_conv.scala 138:36]
  wire  _GEN_8; // @[mmu_conv.scala 133:21]
  wire  _GEN_9; // @[mmu_conv.scala 128:42]
  wire  protect_exception_0; // @[mmu_conv.scala 125:18]
  wire  _GEN_11; // @[mmu_conv.scala 145:32]
  wire  _T_28; // @[mmu_conv.scala 148:36]
  wire  update_exception_0; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_29; // @[Cat.scala 29:58]
  wire [33:0] _GEN_286; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_30; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_32; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_287; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_36; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_37; // @[mmu_conv.scala 113:64]
  wire  _T_38; // @[mmu_conv.scala 113:48]
  wire  _GEN_13; // @[mmu_conv.scala 112:50]
  wire  _GEN_14; // @[mmu_conv.scala 109:45]
  wire  hit_1; // @[mmu_conv.scala 119:32]
  wire  _GEN_16; // @[mmu_conv.scala 126:35]
  wire  _GEN_17; // @[mmu_conv.scala 129:35]
  wire  _GEN_18; // @[mmu_conv.scala 130:35]
  wire  _T_53; // @[mmu_conv.scala 134:36]
  wire  _GEN_19; // @[mmu_conv.scala 134:61]
  wire  _GEN_20; // @[mmu_conv.scala 138:36]
  wire  _GEN_21; // @[mmu_conv.scala 133:21]
  wire  _GEN_22; // @[mmu_conv.scala 128:42]
  wire  protect_exception_1; // @[mmu_conv.scala 125:18]
  wire  _GEN_24; // @[mmu_conv.scala 145:32]
  wire  _T_62; // @[mmu_conv.scala 148:36]
  wire  update_exception_1; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_63; // @[Cat.scala 29:58]
  wire [33:0] _GEN_288; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_64; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_66; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_289; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_70; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_71; // @[mmu_conv.scala 113:64]
  wire  _T_72; // @[mmu_conv.scala 113:48]
  wire  _GEN_26; // @[mmu_conv.scala 112:50]
  wire  _GEN_27; // @[mmu_conv.scala 109:45]
  wire  hit_2; // @[mmu_conv.scala 119:32]
  wire  _GEN_29; // @[mmu_conv.scala 126:35]
  wire  _GEN_30; // @[mmu_conv.scala 129:35]
  wire  _GEN_31; // @[mmu_conv.scala 130:35]
  wire  _T_87; // @[mmu_conv.scala 134:36]
  wire  _GEN_32; // @[mmu_conv.scala 134:61]
  wire  _GEN_33; // @[mmu_conv.scala 138:36]
  wire  _GEN_34; // @[mmu_conv.scala 133:21]
  wire  _GEN_35; // @[mmu_conv.scala 128:42]
  wire  protect_exception_2; // @[mmu_conv.scala 125:18]
  wire  _GEN_37; // @[mmu_conv.scala 145:32]
  wire  _T_96; // @[mmu_conv.scala 148:36]
  wire  update_exception_2; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_97; // @[Cat.scala 29:58]
  wire [33:0] _GEN_290; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_98; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_100; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_291; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_104; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_105; // @[mmu_conv.scala 113:64]
  wire  _T_106; // @[mmu_conv.scala 113:48]
  wire  _GEN_39; // @[mmu_conv.scala 112:50]
  wire  _GEN_40; // @[mmu_conv.scala 109:45]
  wire  hit_3; // @[mmu_conv.scala 119:32]
  wire  _GEN_42; // @[mmu_conv.scala 126:35]
  wire  _GEN_43; // @[mmu_conv.scala 129:35]
  wire  _GEN_44; // @[mmu_conv.scala 130:35]
  wire  _T_121; // @[mmu_conv.scala 134:36]
  wire  _GEN_45; // @[mmu_conv.scala 134:61]
  wire  _GEN_46; // @[mmu_conv.scala 138:36]
  wire  _GEN_47; // @[mmu_conv.scala 133:21]
  wire  _GEN_48; // @[mmu_conv.scala 128:42]
  wire  protect_exception_3; // @[mmu_conv.scala 125:18]
  wire  _GEN_50; // @[mmu_conv.scala 145:32]
  wire  _T_130; // @[mmu_conv.scala 148:36]
  wire  update_exception_3; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_131; // @[Cat.scala 29:58]
  wire [33:0] _GEN_292; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_132; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_134; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_293; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_138; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_139; // @[mmu_conv.scala 113:64]
  wire  _T_140; // @[mmu_conv.scala 113:48]
  wire  _GEN_52; // @[mmu_conv.scala 112:50]
  wire  _GEN_53; // @[mmu_conv.scala 109:45]
  wire  hit_4; // @[mmu_conv.scala 119:32]
  wire  _GEN_55; // @[mmu_conv.scala 126:35]
  wire  _GEN_56; // @[mmu_conv.scala 129:35]
  wire  _GEN_57; // @[mmu_conv.scala 130:35]
  wire  _T_155; // @[mmu_conv.scala 134:36]
  wire  _GEN_58; // @[mmu_conv.scala 134:61]
  wire  _GEN_59; // @[mmu_conv.scala 138:36]
  wire  _GEN_60; // @[mmu_conv.scala 133:21]
  wire  _GEN_61; // @[mmu_conv.scala 128:42]
  wire  protect_exception_4; // @[mmu_conv.scala 125:18]
  wire  _GEN_63; // @[mmu_conv.scala 145:32]
  wire  _T_164; // @[mmu_conv.scala 148:36]
  wire  update_exception_4; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_165; // @[Cat.scala 29:58]
  wire [33:0] _GEN_294; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_166; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_168; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_295; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_172; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_173; // @[mmu_conv.scala 113:64]
  wire  _T_174; // @[mmu_conv.scala 113:48]
  wire  _GEN_65; // @[mmu_conv.scala 112:50]
  wire  _GEN_66; // @[mmu_conv.scala 109:45]
  wire  hit_5; // @[mmu_conv.scala 119:32]
  wire  _GEN_68; // @[mmu_conv.scala 126:35]
  wire  _GEN_69; // @[mmu_conv.scala 129:35]
  wire  _GEN_70; // @[mmu_conv.scala 130:35]
  wire  _T_189; // @[mmu_conv.scala 134:36]
  wire  _GEN_71; // @[mmu_conv.scala 134:61]
  wire  _GEN_72; // @[mmu_conv.scala 138:36]
  wire  _GEN_73; // @[mmu_conv.scala 133:21]
  wire  _GEN_74; // @[mmu_conv.scala 128:42]
  wire  protect_exception_5; // @[mmu_conv.scala 125:18]
  wire  _GEN_76; // @[mmu_conv.scala 145:32]
  wire  _T_198; // @[mmu_conv.scala 148:36]
  wire  update_exception_5; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_199; // @[Cat.scala 29:58]
  wire [33:0] _GEN_296; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_200; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_202; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_297; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_206; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_207; // @[mmu_conv.scala 113:64]
  wire  _T_208; // @[mmu_conv.scala 113:48]
  wire  _GEN_78; // @[mmu_conv.scala 112:50]
  wire  _GEN_79; // @[mmu_conv.scala 109:45]
  wire  hit_6; // @[mmu_conv.scala 119:32]
  wire  _GEN_81; // @[mmu_conv.scala 126:35]
  wire  _GEN_82; // @[mmu_conv.scala 129:35]
  wire  _GEN_83; // @[mmu_conv.scala 130:35]
  wire  _T_223; // @[mmu_conv.scala 134:36]
  wire  _GEN_84; // @[mmu_conv.scala 134:61]
  wire  _GEN_85; // @[mmu_conv.scala 138:36]
  wire  _GEN_86; // @[mmu_conv.scala 133:21]
  wire  _GEN_87; // @[mmu_conv.scala 128:42]
  wire  protect_exception_6; // @[mmu_conv.scala 125:18]
  wire  _GEN_89; // @[mmu_conv.scala 145:32]
  wire  _T_232; // @[mmu_conv.scala 148:36]
  wire  update_exception_6; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_233; // @[Cat.scala 29:58]
  wire [33:0] _GEN_298; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_234; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_236; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_299; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_240; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_241; // @[mmu_conv.scala 113:64]
  wire  _T_242; // @[mmu_conv.scala 113:48]
  wire  _GEN_91; // @[mmu_conv.scala 112:50]
  wire  _GEN_92; // @[mmu_conv.scala 109:45]
  wire  hit_7; // @[mmu_conv.scala 119:32]
  wire  _GEN_94; // @[mmu_conv.scala 126:35]
  wire  _GEN_95; // @[mmu_conv.scala 129:35]
  wire  _GEN_96; // @[mmu_conv.scala 130:35]
  wire  _T_257; // @[mmu_conv.scala 134:36]
  wire  _GEN_97; // @[mmu_conv.scala 134:61]
  wire  _GEN_98; // @[mmu_conv.scala 138:36]
  wire  _GEN_99; // @[mmu_conv.scala 133:21]
  wire  _GEN_100; // @[mmu_conv.scala 128:42]
  wire  protect_exception_7; // @[mmu_conv.scala 125:18]
  wire  _GEN_102; // @[mmu_conv.scala 145:32]
  wire  _T_266; // @[mmu_conv.scala 148:36]
  wire  update_exception_7; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_267; // @[Cat.scala 29:58]
  wire [33:0] _GEN_300; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_268; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_270; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_301; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_274; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_275; // @[mmu_conv.scala 113:64]
  wire  _T_276; // @[mmu_conv.scala 113:48]
  wire  _GEN_104; // @[mmu_conv.scala 112:50]
  wire  _GEN_105; // @[mmu_conv.scala 109:45]
  wire  hit_8; // @[mmu_conv.scala 119:32]
  wire  _GEN_107; // @[mmu_conv.scala 126:35]
  wire  _GEN_108; // @[mmu_conv.scala 129:35]
  wire  _GEN_109; // @[mmu_conv.scala 130:35]
  wire  _T_291; // @[mmu_conv.scala 134:36]
  wire  _GEN_110; // @[mmu_conv.scala 134:61]
  wire  _GEN_111; // @[mmu_conv.scala 138:36]
  wire  _GEN_112; // @[mmu_conv.scala 133:21]
  wire  _GEN_113; // @[mmu_conv.scala 128:42]
  wire  protect_exception_8; // @[mmu_conv.scala 125:18]
  wire  _GEN_115; // @[mmu_conv.scala 145:32]
  wire  _T_300; // @[mmu_conv.scala 148:36]
  wire  update_exception_8; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_301; // @[Cat.scala 29:58]
  wire [33:0] _GEN_302; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_302; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_304; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_303; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_308; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_309; // @[mmu_conv.scala 113:64]
  wire  _T_310; // @[mmu_conv.scala 113:48]
  wire  _GEN_117; // @[mmu_conv.scala 112:50]
  wire  _GEN_118; // @[mmu_conv.scala 109:45]
  wire  hit_9; // @[mmu_conv.scala 119:32]
  wire  _GEN_120; // @[mmu_conv.scala 126:35]
  wire  _GEN_121; // @[mmu_conv.scala 129:35]
  wire  _GEN_122; // @[mmu_conv.scala 130:35]
  wire  _T_325; // @[mmu_conv.scala 134:36]
  wire  _GEN_123; // @[mmu_conv.scala 134:61]
  wire  _GEN_124; // @[mmu_conv.scala 138:36]
  wire  _GEN_125; // @[mmu_conv.scala 133:21]
  wire  _GEN_126; // @[mmu_conv.scala 128:42]
  wire  protect_exception_9; // @[mmu_conv.scala 125:18]
  wire  _GEN_128; // @[mmu_conv.scala 145:32]
  wire  _T_334; // @[mmu_conv.scala 148:36]
  wire  update_exception_9; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_335; // @[Cat.scala 29:58]
  wire [33:0] _GEN_304; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_336; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_338; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_305; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_342; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_343; // @[mmu_conv.scala 113:64]
  wire  _T_344; // @[mmu_conv.scala 113:48]
  wire  _GEN_130; // @[mmu_conv.scala 112:50]
  wire  _GEN_131; // @[mmu_conv.scala 109:45]
  wire  hit_10; // @[mmu_conv.scala 119:32]
  wire  _GEN_133; // @[mmu_conv.scala 126:35]
  wire  _GEN_134; // @[mmu_conv.scala 129:35]
  wire  _GEN_135; // @[mmu_conv.scala 130:35]
  wire  _T_359; // @[mmu_conv.scala 134:36]
  wire  _GEN_136; // @[mmu_conv.scala 134:61]
  wire  _GEN_137; // @[mmu_conv.scala 138:36]
  wire  _GEN_138; // @[mmu_conv.scala 133:21]
  wire  _GEN_139; // @[mmu_conv.scala 128:42]
  wire  protect_exception_10; // @[mmu_conv.scala 125:18]
  wire  _GEN_141; // @[mmu_conv.scala 145:32]
  wire  _T_368; // @[mmu_conv.scala 148:36]
  wire  update_exception_10; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_369; // @[Cat.scala 29:58]
  wire [33:0] _GEN_306; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_370; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_372; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_307; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_376; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_377; // @[mmu_conv.scala 113:64]
  wire  _T_378; // @[mmu_conv.scala 113:48]
  wire  _GEN_143; // @[mmu_conv.scala 112:50]
  wire  _GEN_144; // @[mmu_conv.scala 109:45]
  wire  hit_11; // @[mmu_conv.scala 119:32]
  wire  _GEN_146; // @[mmu_conv.scala 126:35]
  wire  _GEN_147; // @[mmu_conv.scala 129:35]
  wire  _GEN_148; // @[mmu_conv.scala 130:35]
  wire  _T_393; // @[mmu_conv.scala 134:36]
  wire  _GEN_149; // @[mmu_conv.scala 134:61]
  wire  _GEN_150; // @[mmu_conv.scala 138:36]
  wire  _GEN_151; // @[mmu_conv.scala 133:21]
  wire  _GEN_152; // @[mmu_conv.scala 128:42]
  wire  protect_exception_11; // @[mmu_conv.scala 125:18]
  wire  _GEN_154; // @[mmu_conv.scala 145:32]
  wire  _T_402; // @[mmu_conv.scala 148:36]
  wire  update_exception_11; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_403; // @[Cat.scala 29:58]
  wire [33:0] _GEN_308; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_404; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_406; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_309; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_410; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_411; // @[mmu_conv.scala 113:64]
  wire  _T_412; // @[mmu_conv.scala 113:48]
  wire  _GEN_156; // @[mmu_conv.scala 112:50]
  wire  _GEN_157; // @[mmu_conv.scala 109:45]
  wire  hit_12; // @[mmu_conv.scala 119:32]
  wire  _GEN_159; // @[mmu_conv.scala 126:35]
  wire  _GEN_160; // @[mmu_conv.scala 129:35]
  wire  _GEN_161; // @[mmu_conv.scala 130:35]
  wire  _T_427; // @[mmu_conv.scala 134:36]
  wire  _GEN_162; // @[mmu_conv.scala 134:61]
  wire  _GEN_163; // @[mmu_conv.scala 138:36]
  wire  _GEN_164; // @[mmu_conv.scala 133:21]
  wire  _GEN_165; // @[mmu_conv.scala 128:42]
  wire  protect_exception_12; // @[mmu_conv.scala 125:18]
  wire  _GEN_167; // @[mmu_conv.scala 145:32]
  wire  _T_436; // @[mmu_conv.scala 148:36]
  wire  update_exception_12; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_437; // @[Cat.scala 29:58]
  wire [33:0] _GEN_310; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_438; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_440; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_311; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_444; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_445; // @[mmu_conv.scala 113:64]
  wire  _T_446; // @[mmu_conv.scala 113:48]
  wire  _GEN_169; // @[mmu_conv.scala 112:50]
  wire  _GEN_170; // @[mmu_conv.scala 109:45]
  wire  hit_13; // @[mmu_conv.scala 119:32]
  wire  _GEN_172; // @[mmu_conv.scala 126:35]
  wire  _GEN_173; // @[mmu_conv.scala 129:35]
  wire  _GEN_174; // @[mmu_conv.scala 130:35]
  wire  _T_461; // @[mmu_conv.scala 134:36]
  wire  _GEN_175; // @[mmu_conv.scala 134:61]
  wire  _GEN_176; // @[mmu_conv.scala 138:36]
  wire  _GEN_177; // @[mmu_conv.scala 133:21]
  wire  _GEN_178; // @[mmu_conv.scala 128:42]
  wire  protect_exception_13; // @[mmu_conv.scala 125:18]
  wire  _GEN_180; // @[mmu_conv.scala 145:32]
  wire  _T_470; // @[mmu_conv.scala 148:36]
  wire  update_exception_13; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_471; // @[Cat.scala 29:58]
  wire [33:0] _GEN_312; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_472; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_474; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_313; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_478; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_479; // @[mmu_conv.scala 113:64]
  wire  _T_480; // @[mmu_conv.scala 113:48]
  wire  _GEN_182; // @[mmu_conv.scala 112:50]
  wire  _GEN_183; // @[mmu_conv.scala 109:45]
  wire  hit_14; // @[mmu_conv.scala 119:32]
  wire  _GEN_185; // @[mmu_conv.scala 126:35]
  wire  _GEN_186; // @[mmu_conv.scala 129:35]
  wire  _GEN_187; // @[mmu_conv.scala 130:35]
  wire  _T_495; // @[mmu_conv.scala 134:36]
  wire  _GEN_188; // @[mmu_conv.scala 134:61]
  wire  _GEN_189; // @[mmu_conv.scala 138:36]
  wire  _GEN_190; // @[mmu_conv.scala 133:21]
  wire  _GEN_191; // @[mmu_conv.scala 128:42]
  wire  protect_exception_14; // @[mmu_conv.scala 125:18]
  wire  _GEN_193; // @[mmu_conv.scala 145:32]
  wire  _T_504; // @[mmu_conv.scala 148:36]
  wire  update_exception_14; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_505; // @[Cat.scala 29:58]
  wire [33:0] _GEN_314; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_506; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_508; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_315; // @[mmu_conv.scala 152:62]
  wire [31:0] _T_512; // @[mmu_conv.scala 113:33]
  wire [31:0] _T_513; // @[mmu_conv.scala 113:64]
  wire  _T_514; // @[mmu_conv.scala 113:48]
  wire  _GEN_195; // @[mmu_conv.scala 112:50]
  wire  _GEN_196; // @[mmu_conv.scala 109:45]
  wire  hit_15; // @[mmu_conv.scala 119:32]
  wire  _GEN_198; // @[mmu_conv.scala 126:35]
  wire  _GEN_199; // @[mmu_conv.scala 129:35]
  wire  _GEN_200; // @[mmu_conv.scala 130:35]
  wire  _T_529; // @[mmu_conv.scala 134:36]
  wire  _GEN_201; // @[mmu_conv.scala 134:61]
  wire  _GEN_202; // @[mmu_conv.scala 138:36]
  wire  _GEN_203; // @[mmu_conv.scala 133:21]
  wire  _GEN_204; // @[mmu_conv.scala 128:42]
  wire  protect_exception_15; // @[mmu_conv.scala 125:18]
  wire  _GEN_206; // @[mmu_conv.scala 145:32]
  wire  _T_538; // @[mmu_conv.scala 148:36]
  wire  update_exception_15; // @[mmu_conv.scala 148:61]
  wire [33:0] _T_539; // @[Cat.scala 29:58]
  wire [33:0] _GEN_316; // @[mmu_conv.scala 152:47]
  wire [33:0] _T_540; // @[mmu_conv.scala 152:47]
  wire [31:0] _T_542; // @[mmu_conv.scala 152:79]
  wire [33:0] _GEN_317; // @[mmu_conv.scala 152:62]
  wire [7:0] _T_550; // @[mmu_conv.scala 158:33]
  wire [15:0] _T_558; // @[mmu_conv.scala 158:33]
  wire  _T_559; // @[mmu_conv.scala 158:40]
  wire  tlb_miss_exception; // @[mmu_conv.scala 158:28]
  wire [3:0] _GEN_208; // @[mmu_conv.scala 161:17]
  wire [3:0] _GEN_209; // @[mmu_conv.scala 162:17]
  wire [3:0] _GEN_210; // @[mmu_conv.scala 163:17]
  wire [3:0] _GEN_211; // @[mmu_conv.scala 164:17]
  wire [3:0] _GEN_212; // @[mmu_conv.scala 165:17]
  wire [3:0] _GEN_213; // @[mmu_conv.scala 166:17]
  wire [3:0] _GEN_214; // @[mmu_conv.scala 167:17]
  wire [3:0] _GEN_215; // @[mmu_conv.scala 168:17]
  wire [3:0] _GEN_216; // @[mmu_conv.scala 169:17]
  wire [3:0] _GEN_217; // @[mmu_conv.scala 170:17]
  wire [3:0] _GEN_218; // @[mmu_conv.scala 171:17]
  wire [3:0] _GEN_219; // @[mmu_conv.scala 172:17]
  wire [3:0] _GEN_220; // @[mmu_conv.scala 173:17]
  wire [3:0] _GEN_221; // @[mmu_conv.scala 174:17]
  wire [3:0] _GEN_222; // @[mmu_conv.scala 175:17]
  wire  _GEN_225; // @[mmu_conv.scala 178:39]
  wire  _GEN_226; // @[mmu_conv.scala 178:39]
  wire  _GEN_227; // @[mmu_conv.scala 178:39]
  wire  _GEN_228; // @[mmu_conv.scala 178:39]
  wire  _GEN_229; // @[mmu_conv.scala 178:39]
  wire  _GEN_230; // @[mmu_conv.scala 178:39]
  wire  _GEN_231; // @[mmu_conv.scala 178:39]
  wire  _GEN_232; // @[mmu_conv.scala 178:39]
  wire  _GEN_233; // @[mmu_conv.scala 178:39]
  wire  _GEN_234; // @[mmu_conv.scala 178:39]
  wire  _GEN_235; // @[mmu_conv.scala 178:39]
  wire  _GEN_236; // @[mmu_conv.scala 178:39]
  wire  _GEN_237; // @[mmu_conv.scala 178:39]
  wire  _GEN_238; // @[mmu_conv.scala 178:39]
  wire  _GEN_239; // @[mmu_conv.scala 178:39]
  wire  _T_562; // @[mmu_conv.scala 178:39]
  wire  _GEN_241; // @[mmu_conv.scala 178:75]
  wire  _GEN_242; // @[mmu_conv.scala 178:75]
  wire  _GEN_243; // @[mmu_conv.scala 178:75]
  wire  _GEN_244; // @[mmu_conv.scala 178:75]
  wire  _GEN_245; // @[mmu_conv.scala 178:75]
  wire  _GEN_246; // @[mmu_conv.scala 178:75]
  wire  _GEN_247; // @[mmu_conv.scala 178:75]
  wire  _GEN_248; // @[mmu_conv.scala 178:75]
  wire  _GEN_249; // @[mmu_conv.scala 178:75]
  wire  _GEN_250; // @[mmu_conv.scala 178:75]
  wire  _GEN_251; // @[mmu_conv.scala 178:75]
  wire  _GEN_252; // @[mmu_conv.scala 178:75]
  wire  _GEN_253; // @[mmu_conv.scala 178:75]
  wire  _GEN_254; // @[mmu_conv.scala 178:75]
  wire  _GEN_255; // @[mmu_conv.scala 178:75]
  wire  tlb_exception; // @[mmu_conv.scala 178:75]
  wire  _T_566; // @[mmu_conv.scala 191:23]
  wire  _T_568; // @[mmu_conv.scala 191:35]
  wire [33:0] _GEN_257; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_258; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_259; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_260; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_261; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_262; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_263; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_264; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_265; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_266; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_267; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_268; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_269; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_270; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_271; // @[mmu_conv.scala 201:21]
  wire [33:0] _GEN_272; // @[mmu_conv.scala 200:36]
  wire  _GEN_273; // @[mmu_conv.scala 204:36]
  wire [33:0] _GEN_274; // @[mmu_conv.scala 198:48]
  wire  _GEN_275; // @[mmu_conv.scala 198:48]
  wire  _GEN_276; // @[mmu_conv.scala 198:48]
  wire [33:0] _GEN_277; // @[mmu_conv.scala 191:73]
  wire  _GEN_278; // @[mmu_conv.scala 191:73]
  wire  _GEN_279; // @[mmu_conv.scala 191:73]
  wire [33:0] _GEN_280; // @[mmu_conv.scala 186:40]
  wire  _GEN_281; // @[mmu_conv.scala 186:40]
  wire  _GEN_282; // @[mmu_conv.scala 186:40]
  assign _T = io_vm_i == 5'h0; // @[mmu_conv.scala 109:18]
  assign _T_1 = io_vm_i == 5'h8; // @[mmu_conv.scala 112:24]
  assign _T_2 = io_vir_addr_i & tlb_mask_0; // @[mmu_conv.scala 113:33]
  assign _T_3 = tlb_vpn_0 & tlb_mask_0; // @[mmu_conv.scala 113:64]
  assign _T_4 = _T_2 == _T_3; // @[mmu_conv.scala 113:48]
  assign _GEN_0 = _T_1 & _T_4; // @[mmu_conv.scala 112:50]
  assign _GEN_1 = _T ? 1'h0 : _GEN_0; // @[mmu_conv.scala 109:45]
  assign hit_0 = tlb_pte_0[0] ? _GEN_1 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_3 = ~tlb_pte_0[3] | ~hit_0; // @[mmu_conv.scala 126:35]
  assign _GEN_4 = ~tlb_pte_0[2] | ~hit_0; // @[mmu_conv.scala 129:35]
  assign _GEN_5 = ~tlb_pte_0[1] | _GEN_4; // @[mmu_conv.scala 130:35]
  assign _T_19 = ~tlb_pte_0[1] & ~tlb_pte_0[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_6 = _T_19 | ~hit_0; // @[mmu_conv.scala 134:61]
  assign _GEN_7 = ~tlb_pte_0[1] | ~hit_0; // @[mmu_conv.scala 138:36]
  assign _GEN_8 = io_mxr_i ? _GEN_6 : _GEN_7; // @[mmu_conv.scala 133:21]
  assign _GEN_9 = io_we_i ? _GEN_5 : _GEN_8; // @[mmu_conv.scala 128:42]
  assign protect_exception_0 = io_ex_i ? _GEN_3 : _GEN_9; // @[mmu_conv.scala 125:18]
  assign _GEN_11 = ~tlb_pte_0[6] | ~hit_0; // @[mmu_conv.scala 145:32]
  assign _T_28 = io_we_i & ~tlb_pte_0[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_0 = _T_28 | _GEN_11; // @[mmu_conv.scala 148:61]
  assign _T_29 = {tlb_pte_0,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_286 = {{2'd0}, tlb_mask_0}; // @[mmu_conv.scala 152:47]
  assign _T_30 = _T_29 & _GEN_286; // @[mmu_conv.scala 152:47]
  assign _T_32 = io_vir_addr_i & ~tlb_mask_0; // @[mmu_conv.scala 152:79]
  assign _GEN_287 = {{2'd0}, _T_32}; // @[mmu_conv.scala 152:62]
  assign _T_36 = io_vir_addr_i & tlb_mask_1; // @[mmu_conv.scala 113:33]
  assign _T_37 = tlb_vpn_1 & tlb_mask_1; // @[mmu_conv.scala 113:64]
  assign _T_38 = _T_36 == _T_37; // @[mmu_conv.scala 113:48]
  assign _GEN_13 = _T_1 & _T_38; // @[mmu_conv.scala 112:50]
  assign _GEN_14 = _T ? 1'h0 : _GEN_13; // @[mmu_conv.scala 109:45]
  assign hit_1 = tlb_pte_1[0] ? _GEN_14 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_16 = ~tlb_pte_1[3] | ~hit_1; // @[mmu_conv.scala 126:35]
  assign _GEN_17 = ~tlb_pte_1[2] | ~hit_1; // @[mmu_conv.scala 129:35]
  assign _GEN_18 = ~tlb_pte_1[1] | _GEN_17; // @[mmu_conv.scala 130:35]
  assign _T_53 = ~tlb_pte_1[1] & ~tlb_pte_1[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_19 = _T_53 | ~hit_1; // @[mmu_conv.scala 134:61]
  assign _GEN_20 = ~tlb_pte_1[1] | ~hit_1; // @[mmu_conv.scala 138:36]
  assign _GEN_21 = io_mxr_i ? _GEN_19 : _GEN_20; // @[mmu_conv.scala 133:21]
  assign _GEN_22 = io_we_i ? _GEN_18 : _GEN_21; // @[mmu_conv.scala 128:42]
  assign protect_exception_1 = io_ex_i ? _GEN_16 : _GEN_22; // @[mmu_conv.scala 125:18]
  assign _GEN_24 = ~tlb_pte_1[6] | ~hit_1; // @[mmu_conv.scala 145:32]
  assign _T_62 = io_we_i & ~tlb_pte_1[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_1 = _T_62 | _GEN_24; // @[mmu_conv.scala 148:61]
  assign _T_63 = {tlb_pte_1,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_288 = {{2'd0}, tlb_mask_1}; // @[mmu_conv.scala 152:47]
  assign _T_64 = _T_63 & _GEN_288; // @[mmu_conv.scala 152:47]
  assign _T_66 = io_vir_addr_i & ~tlb_mask_1; // @[mmu_conv.scala 152:79]
  assign _GEN_289 = {{2'd0}, _T_66}; // @[mmu_conv.scala 152:62]
  assign _T_70 = io_vir_addr_i & tlb_mask_2; // @[mmu_conv.scala 113:33]
  assign _T_71 = tlb_vpn_2 & tlb_mask_2; // @[mmu_conv.scala 113:64]
  assign _T_72 = _T_70 == _T_71; // @[mmu_conv.scala 113:48]
  assign _GEN_26 = _T_1 & _T_72; // @[mmu_conv.scala 112:50]
  assign _GEN_27 = _T ? 1'h0 : _GEN_26; // @[mmu_conv.scala 109:45]
  assign hit_2 = tlb_pte_2[0] ? _GEN_27 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_29 = ~tlb_pte_2[3] | ~hit_2; // @[mmu_conv.scala 126:35]
  assign _GEN_30 = ~tlb_pte_2[2] | ~hit_2; // @[mmu_conv.scala 129:35]
  assign _GEN_31 = ~tlb_pte_2[1] | _GEN_30; // @[mmu_conv.scala 130:35]
  assign _T_87 = ~tlb_pte_2[1] & ~tlb_pte_2[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_32 = _T_87 | ~hit_2; // @[mmu_conv.scala 134:61]
  assign _GEN_33 = ~tlb_pte_2[1] | ~hit_2; // @[mmu_conv.scala 138:36]
  assign _GEN_34 = io_mxr_i ? _GEN_32 : _GEN_33; // @[mmu_conv.scala 133:21]
  assign _GEN_35 = io_we_i ? _GEN_31 : _GEN_34; // @[mmu_conv.scala 128:42]
  assign protect_exception_2 = io_ex_i ? _GEN_29 : _GEN_35; // @[mmu_conv.scala 125:18]
  assign _GEN_37 = ~tlb_pte_2[6] | ~hit_2; // @[mmu_conv.scala 145:32]
  assign _T_96 = io_we_i & ~tlb_pte_2[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_2 = _T_96 | _GEN_37; // @[mmu_conv.scala 148:61]
  assign _T_97 = {tlb_pte_2,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_290 = {{2'd0}, tlb_mask_2}; // @[mmu_conv.scala 152:47]
  assign _T_98 = _T_97 & _GEN_290; // @[mmu_conv.scala 152:47]
  assign _T_100 = io_vir_addr_i & ~tlb_mask_2; // @[mmu_conv.scala 152:79]
  assign _GEN_291 = {{2'd0}, _T_100}; // @[mmu_conv.scala 152:62]
  assign _T_104 = io_vir_addr_i & tlb_mask_3; // @[mmu_conv.scala 113:33]
  assign _T_105 = tlb_vpn_3 & tlb_mask_3; // @[mmu_conv.scala 113:64]
  assign _T_106 = _T_104 == _T_105; // @[mmu_conv.scala 113:48]
  assign _GEN_39 = _T_1 & _T_106; // @[mmu_conv.scala 112:50]
  assign _GEN_40 = _T ? 1'h0 : _GEN_39; // @[mmu_conv.scala 109:45]
  assign hit_3 = tlb_pte_3[0] ? _GEN_40 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_42 = ~tlb_pte_3[3] | ~hit_3; // @[mmu_conv.scala 126:35]
  assign _GEN_43 = ~tlb_pte_3[2] | ~hit_3; // @[mmu_conv.scala 129:35]
  assign _GEN_44 = ~tlb_pte_3[1] | _GEN_43; // @[mmu_conv.scala 130:35]
  assign _T_121 = ~tlb_pte_3[1] & ~tlb_pte_3[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_45 = _T_121 | ~hit_3; // @[mmu_conv.scala 134:61]
  assign _GEN_46 = ~tlb_pte_3[1] | ~hit_3; // @[mmu_conv.scala 138:36]
  assign _GEN_47 = io_mxr_i ? _GEN_45 : _GEN_46; // @[mmu_conv.scala 133:21]
  assign _GEN_48 = io_we_i ? _GEN_44 : _GEN_47; // @[mmu_conv.scala 128:42]
  assign protect_exception_3 = io_ex_i ? _GEN_42 : _GEN_48; // @[mmu_conv.scala 125:18]
  assign _GEN_50 = ~tlb_pte_3[6] | ~hit_3; // @[mmu_conv.scala 145:32]
  assign _T_130 = io_we_i & ~tlb_pte_3[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_3 = _T_130 | _GEN_50; // @[mmu_conv.scala 148:61]
  assign _T_131 = {tlb_pte_3,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_292 = {{2'd0}, tlb_mask_3}; // @[mmu_conv.scala 152:47]
  assign _T_132 = _T_131 & _GEN_292; // @[mmu_conv.scala 152:47]
  assign _T_134 = io_vir_addr_i & ~tlb_mask_3; // @[mmu_conv.scala 152:79]
  assign _GEN_293 = {{2'd0}, _T_134}; // @[mmu_conv.scala 152:62]
  assign _T_138 = io_vir_addr_i & tlb_mask_4; // @[mmu_conv.scala 113:33]
  assign _T_139 = tlb_vpn_4 & tlb_mask_4; // @[mmu_conv.scala 113:64]
  assign _T_140 = _T_138 == _T_139; // @[mmu_conv.scala 113:48]
  assign _GEN_52 = _T_1 & _T_140; // @[mmu_conv.scala 112:50]
  assign _GEN_53 = _T ? 1'h0 : _GEN_52; // @[mmu_conv.scala 109:45]
  assign hit_4 = tlb_pte_4[0] ? _GEN_53 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_55 = ~tlb_pte_4[3] | ~hit_4; // @[mmu_conv.scala 126:35]
  assign _GEN_56 = ~tlb_pte_4[2] | ~hit_4; // @[mmu_conv.scala 129:35]
  assign _GEN_57 = ~tlb_pte_4[1] | _GEN_56; // @[mmu_conv.scala 130:35]
  assign _T_155 = ~tlb_pte_4[1] & ~tlb_pte_4[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_58 = _T_155 | ~hit_4; // @[mmu_conv.scala 134:61]
  assign _GEN_59 = ~tlb_pte_4[1] | ~hit_4; // @[mmu_conv.scala 138:36]
  assign _GEN_60 = io_mxr_i ? _GEN_58 : _GEN_59; // @[mmu_conv.scala 133:21]
  assign _GEN_61 = io_we_i ? _GEN_57 : _GEN_60; // @[mmu_conv.scala 128:42]
  assign protect_exception_4 = io_ex_i ? _GEN_55 : _GEN_61; // @[mmu_conv.scala 125:18]
  assign _GEN_63 = ~tlb_pte_4[6] | ~hit_4; // @[mmu_conv.scala 145:32]
  assign _T_164 = io_we_i & ~tlb_pte_4[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_4 = _T_164 | _GEN_63; // @[mmu_conv.scala 148:61]
  assign _T_165 = {tlb_pte_4,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_294 = {{2'd0}, tlb_mask_4}; // @[mmu_conv.scala 152:47]
  assign _T_166 = _T_165 & _GEN_294; // @[mmu_conv.scala 152:47]
  assign _T_168 = io_vir_addr_i & ~tlb_mask_4; // @[mmu_conv.scala 152:79]
  assign _GEN_295 = {{2'd0}, _T_168}; // @[mmu_conv.scala 152:62]
  assign _T_172 = io_vir_addr_i & tlb_mask_5; // @[mmu_conv.scala 113:33]
  assign _T_173 = tlb_vpn_5 & tlb_mask_5; // @[mmu_conv.scala 113:64]
  assign _T_174 = _T_172 == _T_173; // @[mmu_conv.scala 113:48]
  assign _GEN_65 = _T_1 & _T_174; // @[mmu_conv.scala 112:50]
  assign _GEN_66 = _T ? 1'h0 : _GEN_65; // @[mmu_conv.scala 109:45]
  assign hit_5 = tlb_pte_5[0] ? _GEN_66 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_68 = ~tlb_pte_5[3] | ~hit_5; // @[mmu_conv.scala 126:35]
  assign _GEN_69 = ~tlb_pte_5[2] | ~hit_5; // @[mmu_conv.scala 129:35]
  assign _GEN_70 = ~tlb_pte_5[1] | _GEN_69; // @[mmu_conv.scala 130:35]
  assign _T_189 = ~tlb_pte_5[1] & ~tlb_pte_5[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_71 = _T_189 | ~hit_5; // @[mmu_conv.scala 134:61]
  assign _GEN_72 = ~tlb_pte_5[1] | ~hit_5; // @[mmu_conv.scala 138:36]
  assign _GEN_73 = io_mxr_i ? _GEN_71 : _GEN_72; // @[mmu_conv.scala 133:21]
  assign _GEN_74 = io_we_i ? _GEN_70 : _GEN_73; // @[mmu_conv.scala 128:42]
  assign protect_exception_5 = io_ex_i ? _GEN_68 : _GEN_74; // @[mmu_conv.scala 125:18]
  assign _GEN_76 = ~tlb_pte_5[6] | ~hit_5; // @[mmu_conv.scala 145:32]
  assign _T_198 = io_we_i & ~tlb_pte_5[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_5 = _T_198 | _GEN_76; // @[mmu_conv.scala 148:61]
  assign _T_199 = {tlb_pte_5,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_296 = {{2'd0}, tlb_mask_5}; // @[mmu_conv.scala 152:47]
  assign _T_200 = _T_199 & _GEN_296; // @[mmu_conv.scala 152:47]
  assign _T_202 = io_vir_addr_i & ~tlb_mask_5; // @[mmu_conv.scala 152:79]
  assign _GEN_297 = {{2'd0}, _T_202}; // @[mmu_conv.scala 152:62]
  assign _T_206 = io_vir_addr_i & tlb_mask_6; // @[mmu_conv.scala 113:33]
  assign _T_207 = tlb_vpn_6 & tlb_mask_6; // @[mmu_conv.scala 113:64]
  assign _T_208 = _T_206 == _T_207; // @[mmu_conv.scala 113:48]
  assign _GEN_78 = _T_1 & _T_208; // @[mmu_conv.scala 112:50]
  assign _GEN_79 = _T ? 1'h0 : _GEN_78; // @[mmu_conv.scala 109:45]
  assign hit_6 = tlb_pte_6[0] ? _GEN_79 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_81 = ~tlb_pte_6[3] | ~hit_6; // @[mmu_conv.scala 126:35]
  assign _GEN_82 = ~tlb_pte_6[2] | ~hit_6; // @[mmu_conv.scala 129:35]
  assign _GEN_83 = ~tlb_pte_6[1] | _GEN_82; // @[mmu_conv.scala 130:35]
  assign _T_223 = ~tlb_pte_6[1] & ~tlb_pte_6[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_84 = _T_223 | ~hit_6; // @[mmu_conv.scala 134:61]
  assign _GEN_85 = ~tlb_pte_6[1] | ~hit_6; // @[mmu_conv.scala 138:36]
  assign _GEN_86 = io_mxr_i ? _GEN_84 : _GEN_85; // @[mmu_conv.scala 133:21]
  assign _GEN_87 = io_we_i ? _GEN_83 : _GEN_86; // @[mmu_conv.scala 128:42]
  assign protect_exception_6 = io_ex_i ? _GEN_81 : _GEN_87; // @[mmu_conv.scala 125:18]
  assign _GEN_89 = ~tlb_pte_6[6] | ~hit_6; // @[mmu_conv.scala 145:32]
  assign _T_232 = io_we_i & ~tlb_pte_6[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_6 = _T_232 | _GEN_89; // @[mmu_conv.scala 148:61]
  assign _T_233 = {tlb_pte_6,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_298 = {{2'd0}, tlb_mask_6}; // @[mmu_conv.scala 152:47]
  assign _T_234 = _T_233 & _GEN_298; // @[mmu_conv.scala 152:47]
  assign _T_236 = io_vir_addr_i & ~tlb_mask_6; // @[mmu_conv.scala 152:79]
  assign _GEN_299 = {{2'd0}, _T_236}; // @[mmu_conv.scala 152:62]
  assign _T_240 = io_vir_addr_i & tlb_mask_7; // @[mmu_conv.scala 113:33]
  assign _T_241 = tlb_vpn_7 & tlb_mask_7; // @[mmu_conv.scala 113:64]
  assign _T_242 = _T_240 == _T_241; // @[mmu_conv.scala 113:48]
  assign _GEN_91 = _T_1 & _T_242; // @[mmu_conv.scala 112:50]
  assign _GEN_92 = _T ? 1'h0 : _GEN_91; // @[mmu_conv.scala 109:45]
  assign hit_7 = tlb_pte_7[0] ? _GEN_92 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_94 = ~tlb_pte_7[3] | ~hit_7; // @[mmu_conv.scala 126:35]
  assign _GEN_95 = ~tlb_pte_7[2] | ~hit_7; // @[mmu_conv.scala 129:35]
  assign _GEN_96 = ~tlb_pte_7[1] | _GEN_95; // @[mmu_conv.scala 130:35]
  assign _T_257 = ~tlb_pte_7[1] & ~tlb_pte_7[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_97 = _T_257 | ~hit_7; // @[mmu_conv.scala 134:61]
  assign _GEN_98 = ~tlb_pte_7[1] | ~hit_7; // @[mmu_conv.scala 138:36]
  assign _GEN_99 = io_mxr_i ? _GEN_97 : _GEN_98; // @[mmu_conv.scala 133:21]
  assign _GEN_100 = io_we_i ? _GEN_96 : _GEN_99; // @[mmu_conv.scala 128:42]
  assign protect_exception_7 = io_ex_i ? _GEN_94 : _GEN_100; // @[mmu_conv.scala 125:18]
  assign _GEN_102 = ~tlb_pte_7[6] | ~hit_7; // @[mmu_conv.scala 145:32]
  assign _T_266 = io_we_i & ~tlb_pte_7[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_7 = _T_266 | _GEN_102; // @[mmu_conv.scala 148:61]
  assign _T_267 = {tlb_pte_7,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_300 = {{2'd0}, tlb_mask_7}; // @[mmu_conv.scala 152:47]
  assign _T_268 = _T_267 & _GEN_300; // @[mmu_conv.scala 152:47]
  assign _T_270 = io_vir_addr_i & ~tlb_mask_7; // @[mmu_conv.scala 152:79]
  assign _GEN_301 = {{2'd0}, _T_270}; // @[mmu_conv.scala 152:62]
  assign _T_274 = io_vir_addr_i & tlb_mask_8; // @[mmu_conv.scala 113:33]
  assign _T_275 = tlb_vpn_8 & tlb_mask_8; // @[mmu_conv.scala 113:64]
  assign _T_276 = _T_274 == _T_275; // @[mmu_conv.scala 113:48]
  assign _GEN_104 = _T_1 & _T_276; // @[mmu_conv.scala 112:50]
  assign _GEN_105 = _T ? 1'h0 : _GEN_104; // @[mmu_conv.scala 109:45]
  assign hit_8 = tlb_pte_8[0] ? _GEN_105 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_107 = ~tlb_pte_8[3] | ~hit_8; // @[mmu_conv.scala 126:35]
  assign _GEN_108 = ~tlb_pte_8[2] | ~hit_8; // @[mmu_conv.scala 129:35]
  assign _GEN_109 = ~tlb_pte_8[1] | _GEN_108; // @[mmu_conv.scala 130:35]
  assign _T_291 = ~tlb_pte_8[1] & ~tlb_pte_8[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_110 = _T_291 | ~hit_8; // @[mmu_conv.scala 134:61]
  assign _GEN_111 = ~tlb_pte_8[1] | ~hit_8; // @[mmu_conv.scala 138:36]
  assign _GEN_112 = io_mxr_i ? _GEN_110 : _GEN_111; // @[mmu_conv.scala 133:21]
  assign _GEN_113 = io_we_i ? _GEN_109 : _GEN_112; // @[mmu_conv.scala 128:42]
  assign protect_exception_8 = io_ex_i ? _GEN_107 : _GEN_113; // @[mmu_conv.scala 125:18]
  assign _GEN_115 = ~tlb_pte_8[6] | ~hit_8; // @[mmu_conv.scala 145:32]
  assign _T_300 = io_we_i & ~tlb_pte_8[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_8 = _T_300 | _GEN_115; // @[mmu_conv.scala 148:61]
  assign _T_301 = {tlb_pte_8,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_302 = {{2'd0}, tlb_mask_8}; // @[mmu_conv.scala 152:47]
  assign _T_302 = _T_301 & _GEN_302; // @[mmu_conv.scala 152:47]
  assign _T_304 = io_vir_addr_i & ~tlb_mask_8; // @[mmu_conv.scala 152:79]
  assign _GEN_303 = {{2'd0}, _T_304}; // @[mmu_conv.scala 152:62]
  assign _T_308 = io_vir_addr_i & tlb_mask_9; // @[mmu_conv.scala 113:33]
  assign _T_309 = tlb_vpn_9 & tlb_mask_9; // @[mmu_conv.scala 113:64]
  assign _T_310 = _T_308 == _T_309; // @[mmu_conv.scala 113:48]
  assign _GEN_117 = _T_1 & _T_310; // @[mmu_conv.scala 112:50]
  assign _GEN_118 = _T ? 1'h0 : _GEN_117; // @[mmu_conv.scala 109:45]
  assign hit_9 = tlb_pte_9[0] ? _GEN_118 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_120 = ~tlb_pte_9[3] | ~hit_9; // @[mmu_conv.scala 126:35]
  assign _GEN_121 = ~tlb_pte_9[2] | ~hit_9; // @[mmu_conv.scala 129:35]
  assign _GEN_122 = ~tlb_pte_9[1] | _GEN_121; // @[mmu_conv.scala 130:35]
  assign _T_325 = ~tlb_pte_9[1] & ~tlb_pte_9[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_123 = _T_325 | ~hit_9; // @[mmu_conv.scala 134:61]
  assign _GEN_124 = ~tlb_pte_9[1] | ~hit_9; // @[mmu_conv.scala 138:36]
  assign _GEN_125 = io_mxr_i ? _GEN_123 : _GEN_124; // @[mmu_conv.scala 133:21]
  assign _GEN_126 = io_we_i ? _GEN_122 : _GEN_125; // @[mmu_conv.scala 128:42]
  assign protect_exception_9 = io_ex_i ? _GEN_120 : _GEN_126; // @[mmu_conv.scala 125:18]
  assign _GEN_128 = ~tlb_pte_9[6] | ~hit_9; // @[mmu_conv.scala 145:32]
  assign _T_334 = io_we_i & ~tlb_pte_9[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_9 = _T_334 | _GEN_128; // @[mmu_conv.scala 148:61]
  assign _T_335 = {tlb_pte_9,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_304 = {{2'd0}, tlb_mask_9}; // @[mmu_conv.scala 152:47]
  assign _T_336 = _T_335 & _GEN_304; // @[mmu_conv.scala 152:47]
  assign _T_338 = io_vir_addr_i & ~tlb_mask_9; // @[mmu_conv.scala 152:79]
  assign _GEN_305 = {{2'd0}, _T_338}; // @[mmu_conv.scala 152:62]
  assign _T_342 = io_vir_addr_i & tlb_mask_10; // @[mmu_conv.scala 113:33]
  assign _T_343 = tlb_vpn_10 & tlb_mask_10; // @[mmu_conv.scala 113:64]
  assign _T_344 = _T_342 == _T_343; // @[mmu_conv.scala 113:48]
  assign _GEN_130 = _T_1 & _T_344; // @[mmu_conv.scala 112:50]
  assign _GEN_131 = _T ? 1'h0 : _GEN_130; // @[mmu_conv.scala 109:45]
  assign hit_10 = tlb_pte_10[0] ? _GEN_131 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_133 = ~tlb_pte_10[3] | ~hit_10; // @[mmu_conv.scala 126:35]
  assign _GEN_134 = ~tlb_pte_10[2] | ~hit_10; // @[mmu_conv.scala 129:35]
  assign _GEN_135 = ~tlb_pte_10[1] | _GEN_134; // @[mmu_conv.scala 130:35]
  assign _T_359 = ~tlb_pte_10[1] & ~tlb_pte_10[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_136 = _T_359 | ~hit_10; // @[mmu_conv.scala 134:61]
  assign _GEN_137 = ~tlb_pte_10[1] | ~hit_10; // @[mmu_conv.scala 138:36]
  assign _GEN_138 = io_mxr_i ? _GEN_136 : _GEN_137; // @[mmu_conv.scala 133:21]
  assign _GEN_139 = io_we_i ? _GEN_135 : _GEN_138; // @[mmu_conv.scala 128:42]
  assign protect_exception_10 = io_ex_i ? _GEN_133 : _GEN_139; // @[mmu_conv.scala 125:18]
  assign _GEN_141 = ~tlb_pte_10[6] | ~hit_10; // @[mmu_conv.scala 145:32]
  assign _T_368 = io_we_i & ~tlb_pte_10[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_10 = _T_368 | _GEN_141; // @[mmu_conv.scala 148:61]
  assign _T_369 = {tlb_pte_10,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_306 = {{2'd0}, tlb_mask_10}; // @[mmu_conv.scala 152:47]
  assign _T_370 = _T_369 & _GEN_306; // @[mmu_conv.scala 152:47]
  assign _T_372 = io_vir_addr_i & ~tlb_mask_10; // @[mmu_conv.scala 152:79]
  assign _GEN_307 = {{2'd0}, _T_372}; // @[mmu_conv.scala 152:62]
  assign _T_376 = io_vir_addr_i & tlb_mask_11; // @[mmu_conv.scala 113:33]
  assign _T_377 = tlb_vpn_11 & tlb_mask_11; // @[mmu_conv.scala 113:64]
  assign _T_378 = _T_376 == _T_377; // @[mmu_conv.scala 113:48]
  assign _GEN_143 = _T_1 & _T_378; // @[mmu_conv.scala 112:50]
  assign _GEN_144 = _T ? 1'h0 : _GEN_143; // @[mmu_conv.scala 109:45]
  assign hit_11 = tlb_pte_11[0] ? _GEN_144 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_146 = ~tlb_pte_11[3] | ~hit_11; // @[mmu_conv.scala 126:35]
  assign _GEN_147 = ~tlb_pte_11[2] | ~hit_11; // @[mmu_conv.scala 129:35]
  assign _GEN_148 = ~tlb_pte_11[1] | _GEN_147; // @[mmu_conv.scala 130:35]
  assign _T_393 = ~tlb_pte_11[1] & ~tlb_pte_11[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_149 = _T_393 | ~hit_11; // @[mmu_conv.scala 134:61]
  assign _GEN_150 = ~tlb_pte_11[1] | ~hit_11; // @[mmu_conv.scala 138:36]
  assign _GEN_151 = io_mxr_i ? _GEN_149 : _GEN_150; // @[mmu_conv.scala 133:21]
  assign _GEN_152 = io_we_i ? _GEN_148 : _GEN_151; // @[mmu_conv.scala 128:42]
  assign protect_exception_11 = io_ex_i ? _GEN_146 : _GEN_152; // @[mmu_conv.scala 125:18]
  assign _GEN_154 = ~tlb_pte_11[6] | ~hit_11; // @[mmu_conv.scala 145:32]
  assign _T_402 = io_we_i & ~tlb_pte_11[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_11 = _T_402 | _GEN_154; // @[mmu_conv.scala 148:61]
  assign _T_403 = {tlb_pte_11,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_308 = {{2'd0}, tlb_mask_11}; // @[mmu_conv.scala 152:47]
  assign _T_404 = _T_403 & _GEN_308; // @[mmu_conv.scala 152:47]
  assign _T_406 = io_vir_addr_i & ~tlb_mask_11; // @[mmu_conv.scala 152:79]
  assign _GEN_309 = {{2'd0}, _T_406}; // @[mmu_conv.scala 152:62]
  assign _T_410 = io_vir_addr_i & tlb_mask_12; // @[mmu_conv.scala 113:33]
  assign _T_411 = tlb_vpn_12 & tlb_mask_12; // @[mmu_conv.scala 113:64]
  assign _T_412 = _T_410 == _T_411; // @[mmu_conv.scala 113:48]
  assign _GEN_156 = _T_1 & _T_412; // @[mmu_conv.scala 112:50]
  assign _GEN_157 = _T ? 1'h0 : _GEN_156; // @[mmu_conv.scala 109:45]
  assign hit_12 = tlb_pte_12[0] ? _GEN_157 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_159 = ~tlb_pte_12[3] | ~hit_12; // @[mmu_conv.scala 126:35]
  assign _GEN_160 = ~tlb_pte_12[2] | ~hit_12; // @[mmu_conv.scala 129:35]
  assign _GEN_161 = ~tlb_pte_12[1] | _GEN_160; // @[mmu_conv.scala 130:35]
  assign _T_427 = ~tlb_pte_12[1] & ~tlb_pte_12[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_162 = _T_427 | ~hit_12; // @[mmu_conv.scala 134:61]
  assign _GEN_163 = ~tlb_pte_12[1] | ~hit_12; // @[mmu_conv.scala 138:36]
  assign _GEN_164 = io_mxr_i ? _GEN_162 : _GEN_163; // @[mmu_conv.scala 133:21]
  assign _GEN_165 = io_we_i ? _GEN_161 : _GEN_164; // @[mmu_conv.scala 128:42]
  assign protect_exception_12 = io_ex_i ? _GEN_159 : _GEN_165; // @[mmu_conv.scala 125:18]
  assign _GEN_167 = ~tlb_pte_12[6] | ~hit_12; // @[mmu_conv.scala 145:32]
  assign _T_436 = io_we_i & ~tlb_pte_12[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_12 = _T_436 | _GEN_167; // @[mmu_conv.scala 148:61]
  assign _T_437 = {tlb_pte_12,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_310 = {{2'd0}, tlb_mask_12}; // @[mmu_conv.scala 152:47]
  assign _T_438 = _T_437 & _GEN_310; // @[mmu_conv.scala 152:47]
  assign _T_440 = io_vir_addr_i & ~tlb_mask_12; // @[mmu_conv.scala 152:79]
  assign _GEN_311 = {{2'd0}, _T_440}; // @[mmu_conv.scala 152:62]
  assign _T_444 = io_vir_addr_i & tlb_mask_13; // @[mmu_conv.scala 113:33]
  assign _T_445 = tlb_vpn_13 & tlb_mask_13; // @[mmu_conv.scala 113:64]
  assign _T_446 = _T_444 == _T_445; // @[mmu_conv.scala 113:48]
  assign _GEN_169 = _T_1 & _T_446; // @[mmu_conv.scala 112:50]
  assign _GEN_170 = _T ? 1'h0 : _GEN_169; // @[mmu_conv.scala 109:45]
  assign hit_13 = tlb_pte_13[0] ? _GEN_170 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_172 = ~tlb_pte_13[3] | ~hit_13; // @[mmu_conv.scala 126:35]
  assign _GEN_173 = ~tlb_pte_13[2] | ~hit_13; // @[mmu_conv.scala 129:35]
  assign _GEN_174 = ~tlb_pte_13[1] | _GEN_173; // @[mmu_conv.scala 130:35]
  assign _T_461 = ~tlb_pte_13[1] & ~tlb_pte_13[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_175 = _T_461 | ~hit_13; // @[mmu_conv.scala 134:61]
  assign _GEN_176 = ~tlb_pte_13[1] | ~hit_13; // @[mmu_conv.scala 138:36]
  assign _GEN_177 = io_mxr_i ? _GEN_175 : _GEN_176; // @[mmu_conv.scala 133:21]
  assign _GEN_178 = io_we_i ? _GEN_174 : _GEN_177; // @[mmu_conv.scala 128:42]
  assign protect_exception_13 = io_ex_i ? _GEN_172 : _GEN_178; // @[mmu_conv.scala 125:18]
  assign _GEN_180 = ~tlb_pte_13[6] | ~hit_13; // @[mmu_conv.scala 145:32]
  assign _T_470 = io_we_i & ~tlb_pte_13[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_13 = _T_470 | _GEN_180; // @[mmu_conv.scala 148:61]
  assign _T_471 = {tlb_pte_13,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_312 = {{2'd0}, tlb_mask_13}; // @[mmu_conv.scala 152:47]
  assign _T_472 = _T_471 & _GEN_312; // @[mmu_conv.scala 152:47]
  assign _T_474 = io_vir_addr_i & ~tlb_mask_13; // @[mmu_conv.scala 152:79]
  assign _GEN_313 = {{2'd0}, _T_474}; // @[mmu_conv.scala 152:62]
  assign _T_478 = io_vir_addr_i & tlb_mask_14; // @[mmu_conv.scala 113:33]
  assign _T_479 = tlb_vpn_14 & tlb_mask_14; // @[mmu_conv.scala 113:64]
  assign _T_480 = _T_478 == _T_479; // @[mmu_conv.scala 113:48]
  assign _GEN_182 = _T_1 & _T_480; // @[mmu_conv.scala 112:50]
  assign _GEN_183 = _T ? 1'h0 : _GEN_182; // @[mmu_conv.scala 109:45]
  assign hit_14 = tlb_pte_14[0] ? _GEN_183 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_185 = ~tlb_pte_14[3] | ~hit_14; // @[mmu_conv.scala 126:35]
  assign _GEN_186 = ~tlb_pte_14[2] | ~hit_14; // @[mmu_conv.scala 129:35]
  assign _GEN_187 = ~tlb_pte_14[1] | _GEN_186; // @[mmu_conv.scala 130:35]
  assign _T_495 = ~tlb_pte_14[1] & ~tlb_pte_14[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_188 = _T_495 | ~hit_14; // @[mmu_conv.scala 134:61]
  assign _GEN_189 = ~tlb_pte_14[1] | ~hit_14; // @[mmu_conv.scala 138:36]
  assign _GEN_190 = io_mxr_i ? _GEN_188 : _GEN_189; // @[mmu_conv.scala 133:21]
  assign _GEN_191 = io_we_i ? _GEN_187 : _GEN_190; // @[mmu_conv.scala 128:42]
  assign protect_exception_14 = io_ex_i ? _GEN_185 : _GEN_191; // @[mmu_conv.scala 125:18]
  assign _GEN_193 = ~tlb_pte_14[6] | ~hit_14; // @[mmu_conv.scala 145:32]
  assign _T_504 = io_we_i & ~tlb_pte_14[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_14 = _T_504 | _GEN_193; // @[mmu_conv.scala 148:61]
  assign _T_505 = {tlb_pte_14,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_314 = {{2'd0}, tlb_mask_14}; // @[mmu_conv.scala 152:47]
  assign _T_506 = _T_505 & _GEN_314; // @[mmu_conv.scala 152:47]
  assign _T_508 = io_vir_addr_i & ~tlb_mask_14; // @[mmu_conv.scala 152:79]
  assign _GEN_315 = {{2'd0}, _T_508}; // @[mmu_conv.scala 152:62]
  assign _T_512 = io_vir_addr_i & tlb_mask_15; // @[mmu_conv.scala 113:33]
  assign _T_513 = tlb_vpn_15 & tlb_mask_15; // @[mmu_conv.scala 113:64]
  assign _T_514 = _T_512 == _T_513; // @[mmu_conv.scala 113:48]
  assign _GEN_195 = _T_1 & _T_514; // @[mmu_conv.scala 112:50]
  assign _GEN_196 = _T ? 1'h0 : _GEN_195; // @[mmu_conv.scala 109:45]
  assign hit_15 = tlb_pte_15[0] ? _GEN_196 : 1'h0; // @[mmu_conv.scala 119:32]
  assign _GEN_198 = ~tlb_pte_15[3] | ~hit_15; // @[mmu_conv.scala 126:35]
  assign _GEN_199 = ~tlb_pte_15[2] | ~hit_15; // @[mmu_conv.scala 129:35]
  assign _GEN_200 = ~tlb_pte_15[1] | _GEN_199; // @[mmu_conv.scala 130:35]
  assign _T_529 = ~tlb_pte_15[1] & ~tlb_pte_15[3]; // @[mmu_conv.scala 134:36]
  assign _GEN_201 = _T_529 | ~hit_15; // @[mmu_conv.scala 134:61]
  assign _GEN_202 = ~tlb_pte_15[1] | ~hit_15; // @[mmu_conv.scala 138:36]
  assign _GEN_203 = io_mxr_i ? _GEN_201 : _GEN_202; // @[mmu_conv.scala 133:21]
  assign _GEN_204 = io_we_i ? _GEN_200 : _GEN_203; // @[mmu_conv.scala 128:42]
  assign protect_exception_15 = io_ex_i ? _GEN_198 : _GEN_204; // @[mmu_conv.scala 125:18]
  assign _GEN_206 = ~tlb_pte_15[6] | ~hit_15; // @[mmu_conv.scala 145:32]
  assign _T_538 = io_we_i & ~tlb_pte_15[7]; // @[mmu_conv.scala 148:36]
  assign update_exception_15 = _T_538 | _GEN_206; // @[mmu_conv.scala 148:61]
  assign _T_539 = {tlb_pte_15,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_316 = {{2'd0}, tlb_mask_15}; // @[mmu_conv.scala 152:47]
  assign _T_540 = _T_539 & _GEN_316; // @[mmu_conv.scala 152:47]
  assign _T_542 = io_vir_addr_i & ~tlb_mask_15; // @[mmu_conv.scala 152:79]
  assign _GEN_317 = {{2'd0}, _T_542}; // @[mmu_conv.scala 152:62]
  assign _T_550 = {hit_7,hit_6,hit_5,hit_4,hit_3,hit_2,hit_1,hit_0}; // @[mmu_conv.scala 158:33]
  assign _T_558 = {hit_15,hit_14,hit_13,hit_12,hit_11,hit_10,hit_9,hit_8,_T_550}; // @[mmu_conv.scala 158:33]
  assign _T_559 = _T_558 != 16'h0; // @[mmu_conv.scala 158:40]
  assign tlb_miss_exception = _T_559 ? 1'h0 : 1'h1; // @[mmu_conv.scala 158:28]
  assign _GEN_208 = hit_15 ? 4'hf : 4'h0; // @[mmu_conv.scala 161:17]
  assign _GEN_209 = hit_14 ? 4'he : _GEN_208; // @[mmu_conv.scala 162:17]
  assign _GEN_210 = hit_13 ? 4'hd : _GEN_209; // @[mmu_conv.scala 163:17]
  assign _GEN_211 = hit_12 ? 4'hc : _GEN_210; // @[mmu_conv.scala 164:17]
  assign _GEN_212 = hit_11 ? 4'hb : _GEN_211; // @[mmu_conv.scala 165:17]
  assign _GEN_213 = hit_10 ? 4'ha : _GEN_212; // @[mmu_conv.scala 166:17]
  assign _GEN_214 = hit_9 ? 4'h9 : _GEN_213; // @[mmu_conv.scala 167:17]
  assign _GEN_215 = hit_8 ? 4'h8 : _GEN_214; // @[mmu_conv.scala 168:17]
  assign _GEN_216 = hit_7 ? 4'h7 : _GEN_215; // @[mmu_conv.scala 169:17]
  assign _GEN_217 = hit_6 ? 4'h6 : _GEN_216; // @[mmu_conv.scala 170:17]
  assign _GEN_218 = hit_5 ? 4'h5 : _GEN_217; // @[mmu_conv.scala 171:17]
  assign _GEN_219 = hit_4 ? 4'h4 : _GEN_218; // @[mmu_conv.scala 172:17]
  assign _GEN_220 = hit_3 ? 4'h3 : _GEN_219; // @[mmu_conv.scala 173:17]
  assign _GEN_221 = hit_2 ? 4'h2 : _GEN_220; // @[mmu_conv.scala 174:17]
  assign _GEN_222 = hit_1 ? 4'h1 : _GEN_221; // @[mmu_conv.scala 175:17]
  assign _GEN_225 = 4'h1 == io_hit_index_o ? protect_exception_1 : protect_exception_0; // @[mmu_conv.scala 178:39]
  assign _GEN_226 = 4'h2 == io_hit_index_o ? protect_exception_2 : _GEN_225; // @[mmu_conv.scala 178:39]
  assign _GEN_227 = 4'h3 == io_hit_index_o ? protect_exception_3 : _GEN_226; // @[mmu_conv.scala 178:39]
  assign _GEN_228 = 4'h4 == io_hit_index_o ? protect_exception_4 : _GEN_227; // @[mmu_conv.scala 178:39]
  assign _GEN_229 = 4'h5 == io_hit_index_o ? protect_exception_5 : _GEN_228; // @[mmu_conv.scala 178:39]
  assign _GEN_230 = 4'h6 == io_hit_index_o ? protect_exception_6 : _GEN_229; // @[mmu_conv.scala 178:39]
  assign _GEN_231 = 4'h7 == io_hit_index_o ? protect_exception_7 : _GEN_230; // @[mmu_conv.scala 178:39]
  assign _GEN_232 = 4'h8 == io_hit_index_o ? protect_exception_8 : _GEN_231; // @[mmu_conv.scala 178:39]
  assign _GEN_233 = 4'h9 == io_hit_index_o ? protect_exception_9 : _GEN_232; // @[mmu_conv.scala 178:39]
  assign _GEN_234 = 4'ha == io_hit_index_o ? protect_exception_10 : _GEN_233; // @[mmu_conv.scala 178:39]
  assign _GEN_235 = 4'hb == io_hit_index_o ? protect_exception_11 : _GEN_234; // @[mmu_conv.scala 178:39]
  assign _GEN_236 = 4'hc == io_hit_index_o ? protect_exception_12 : _GEN_235; // @[mmu_conv.scala 178:39]
  assign _GEN_237 = 4'hd == io_hit_index_o ? protect_exception_13 : _GEN_236; // @[mmu_conv.scala 178:39]
  assign _GEN_238 = 4'he == io_hit_index_o ? protect_exception_14 : _GEN_237; // @[mmu_conv.scala 178:39]
  assign _GEN_239 = 4'hf == io_hit_index_o ? protect_exception_15 : _GEN_238; // @[mmu_conv.scala 178:39]
  assign _T_562 = tlb_miss_exception | _GEN_239; // @[mmu_conv.scala 178:39]
  assign _GEN_241 = 4'h1 == io_hit_index_o ? update_exception_1 : update_exception_0; // @[mmu_conv.scala 178:75]
  assign _GEN_242 = 4'h2 == io_hit_index_o ? update_exception_2 : _GEN_241; // @[mmu_conv.scala 178:75]
  assign _GEN_243 = 4'h3 == io_hit_index_o ? update_exception_3 : _GEN_242; // @[mmu_conv.scala 178:75]
  assign _GEN_244 = 4'h4 == io_hit_index_o ? update_exception_4 : _GEN_243; // @[mmu_conv.scala 178:75]
  assign _GEN_245 = 4'h5 == io_hit_index_o ? update_exception_5 : _GEN_244; // @[mmu_conv.scala 178:75]
  assign _GEN_246 = 4'h6 == io_hit_index_o ? update_exception_6 : _GEN_245; // @[mmu_conv.scala 178:75]
  assign _GEN_247 = 4'h7 == io_hit_index_o ? update_exception_7 : _GEN_246; // @[mmu_conv.scala 178:75]
  assign _GEN_248 = 4'h8 == io_hit_index_o ? update_exception_8 : _GEN_247; // @[mmu_conv.scala 178:75]
  assign _GEN_249 = 4'h9 == io_hit_index_o ? update_exception_9 : _GEN_248; // @[mmu_conv.scala 178:75]
  assign _GEN_250 = 4'ha == io_hit_index_o ? update_exception_10 : _GEN_249; // @[mmu_conv.scala 178:75]
  assign _GEN_251 = 4'hb == io_hit_index_o ? update_exception_11 : _GEN_250; // @[mmu_conv.scala 178:75]
  assign _GEN_252 = 4'hc == io_hit_index_o ? update_exception_12 : _GEN_251; // @[mmu_conv.scala 178:75]
  assign _GEN_253 = 4'hd == io_hit_index_o ? update_exception_13 : _GEN_252; // @[mmu_conv.scala 178:75]
  assign _GEN_254 = 4'he == io_hit_index_o ? update_exception_14 : _GEN_253; // @[mmu_conv.scala 178:75]
  assign _GEN_255 = 4'hf == io_hit_index_o ? update_exception_15 : _GEN_254; // @[mmu_conv.scala 178:75]
  assign tlb_exception = _T_562 | _GEN_255; // @[mmu_conv.scala 178:75]
  assign _T_566 = io_prv_i == 2'h3; // @[mmu_conv.scala 191:23]
  assign _T_568 = _T_566 | _T; // @[mmu_conv.scala 191:35]
  assign _GEN_257 = 4'h1 == io_hit_index_o ? phy_addr_1 : phy_addr_0; // @[mmu_conv.scala 201:21]
  assign _GEN_258 = 4'h2 == io_hit_index_o ? phy_addr_2 : _GEN_257; // @[mmu_conv.scala 201:21]
  assign _GEN_259 = 4'h3 == io_hit_index_o ? phy_addr_3 : _GEN_258; // @[mmu_conv.scala 201:21]
  assign _GEN_260 = 4'h4 == io_hit_index_o ? phy_addr_4 : _GEN_259; // @[mmu_conv.scala 201:21]
  assign _GEN_261 = 4'h5 == io_hit_index_o ? phy_addr_5 : _GEN_260; // @[mmu_conv.scala 201:21]
  assign _GEN_262 = 4'h6 == io_hit_index_o ? phy_addr_6 : _GEN_261; // @[mmu_conv.scala 201:21]
  assign _GEN_263 = 4'h7 == io_hit_index_o ? phy_addr_7 : _GEN_262; // @[mmu_conv.scala 201:21]
  assign _GEN_264 = 4'h8 == io_hit_index_o ? phy_addr_8 : _GEN_263; // @[mmu_conv.scala 201:21]
  assign _GEN_265 = 4'h9 == io_hit_index_o ? phy_addr_9 : _GEN_264; // @[mmu_conv.scala 201:21]
  assign _GEN_266 = 4'ha == io_hit_index_o ? phy_addr_10 : _GEN_265; // @[mmu_conv.scala 201:21]
  assign _GEN_267 = 4'hb == io_hit_index_o ? phy_addr_11 : _GEN_266; // @[mmu_conv.scala 201:21]
  assign _GEN_268 = 4'hc == io_hit_index_o ? phy_addr_12 : _GEN_267; // @[mmu_conv.scala 201:21]
  assign _GEN_269 = 4'hd == io_hit_index_o ? phy_addr_13 : _GEN_268; // @[mmu_conv.scala 201:21]
  assign _GEN_270 = 4'he == io_hit_index_o ? phy_addr_14 : _GEN_269; // @[mmu_conv.scala 201:21]
  assign _GEN_271 = 4'hf == io_hit_index_o ? phy_addr_15 : _GEN_270; // @[mmu_conv.scala 201:21]
  assign _GEN_272 = tlb_exception ? 34'h0 : _GEN_271; // @[mmu_conv.scala 200:36]
  assign _GEN_273 = tlb_miss_exception ? 1'h0 : _GEN_255; // @[mmu_conv.scala 204:36]
  assign _GEN_274 = _T_1 ? _GEN_272 : 34'h0; // @[mmu_conv.scala 198:48]
  assign _GEN_275 = _T_1 & tlb_exception; // @[mmu_conv.scala 198:48]
  assign _GEN_276 = _T_1 & _GEN_273; // @[mmu_conv.scala 198:48]
  assign _GEN_277 = _T_568 ? {{2'd0}, io_vir_addr_i} : _GEN_274; // @[mmu_conv.scala 191:73]
  assign _GEN_278 = _T_568 ? 1'h0 : _GEN_275; // @[mmu_conv.scala 191:73]
  assign _GEN_279 = _T_568 ? 1'h0 : _GEN_276; // @[mmu_conv.scala 191:73]
  assign _GEN_280 = io_ce_i ? _GEN_277 : 34'h0; // @[mmu_conv.scala 186:40]
  assign _GEN_281 = io_ce_i ? _GEN_278 : 1'h0; // @[mmu_conv.scala 186:40]
  assign _GEN_282 = io_ce_i ? _GEN_279 : 1'h0; // @[mmu_conv.scala 186:40]
  assign io_phy_addr_o = io_rst_n ? _GEN_280 : 34'h0; // @[mmu_conv.scala 182:19 mmu_conv.scala 187:19 mmu_conv.scala 192:19 mmu_conv.scala 193:19 mmu_conv.scala 199:19 mmu_conv.scala 201:21 mmu_conv.scala 211:19]
  assign io_tlb_exception_o = io_rst_n ? _GEN_281 : 1'h0; // @[mmu_conv.scala 183:24 mmu_conv.scala 188:24 mmu_conv.scala 195:24 mmu_conv.scala 203:24 mmu_conv.scala 212:24]
  assign io_tlb_update_o = io_rst_n ? _GEN_282 : 1'h0; // @[mmu_conv.scala 184:21 mmu_conv.scala 189:21 mmu_conv.scala 196:21 mmu_conv.scala 205:23 mmu_conv.scala 207:23 mmu_conv.scala 213:21]
  assign io_hit_index_o = hit_0 ? 4'h0 : _GEN_222; // @[mmu_conv.scala 160:18 mmu_conv.scala 161:33 mmu_conv.scala 162:33 mmu_conv.scala 163:33 mmu_conv.scala 164:33 mmu_conv.scala 165:33 mmu_conv.scala 166:33 mmu_conv.scala 167:33 mmu_conv.scala 168:33 mmu_conv.scala 169:33 mmu_conv.scala 170:33 mmu_conv.scala 171:33 mmu_conv.scala 172:33 mmu_conv.scala 173:33 mmu_conv.scala 174:33 mmu_conv.scala 175:33 mmu_conv.scala 176:33]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  tlb_vpn_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tlb_vpn_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  tlb_vpn_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  tlb_vpn_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  tlb_vpn_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  tlb_vpn_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  tlb_vpn_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  tlb_vpn_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  tlb_vpn_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  tlb_vpn_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  tlb_vpn_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  tlb_vpn_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  tlb_vpn_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  tlb_vpn_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  tlb_vpn_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  tlb_vpn_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  tlb_pte_0 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  tlb_pte_1 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  tlb_pte_2 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  tlb_pte_3 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  tlb_pte_4 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  tlb_pte_5 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  tlb_pte_6 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  tlb_pte_7 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  tlb_pte_8 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  tlb_pte_9 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  tlb_pte_10 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  tlb_pte_11 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  tlb_pte_12 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  tlb_pte_13 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  tlb_pte_14 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  tlb_pte_15 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  tlb_mask_0 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  tlb_mask_1 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  tlb_mask_2 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  tlb_mask_3 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  tlb_mask_4 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  tlb_mask_5 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  tlb_mask_6 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  tlb_mask_7 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  tlb_mask_8 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  tlb_mask_9 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  tlb_mask_10 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  tlb_mask_11 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  tlb_mask_12 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  tlb_mask_13 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  tlb_mask_14 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  tlb_mask_15 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {2{`RANDOM}};
  phy_addr_0 = _RAND_48[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {2{`RANDOM}};
  phy_addr_1 = _RAND_49[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {2{`RANDOM}};
  phy_addr_2 = _RAND_50[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {2{`RANDOM}};
  phy_addr_3 = _RAND_51[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {2{`RANDOM}};
  phy_addr_4 = _RAND_52[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {2{`RANDOM}};
  phy_addr_5 = _RAND_53[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {2{`RANDOM}};
  phy_addr_6 = _RAND_54[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {2{`RANDOM}};
  phy_addr_7 = _RAND_55[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {2{`RANDOM}};
  phy_addr_8 = _RAND_56[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {2{`RANDOM}};
  phy_addr_9 = _RAND_57[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {2{`RANDOM}};
  phy_addr_10 = _RAND_58[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {2{`RANDOM}};
  phy_addr_11 = _RAND_59[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {2{`RANDOM}};
  phy_addr_12 = _RAND_60[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {2{`RANDOM}};
  phy_addr_13 = _RAND_61[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {2{`RANDOM}};
  phy_addr_14 = _RAND_62[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {2{`RANDOM}};
  phy_addr_15 = _RAND_63[33:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(*) begin
    tlb_vpn_0 <= io_tlb0_vpn_i;
    tlb_vpn_1 <= io_tlb1_vpn_i;
    tlb_vpn_2 <= io_tlb2_vpn_i;
    tlb_vpn_3 <= io_tlb3_vpn_i;
    tlb_vpn_4 <= io_tlb4_vpn_i;
    tlb_vpn_5 <= io_tlb5_vpn_i;
    tlb_vpn_6 <= io_tlb6_vpn_i;
    tlb_vpn_7 <= io_tlb7_vpn_i;
    tlb_vpn_8 <= io_tlb8_vpn_i;
    tlb_vpn_9 <= io_tlb9_vpn_i;
    tlb_vpn_10 <= io_tlb10_vpn_i;
    tlb_vpn_11 <= io_tlb11_vpn_i;
    tlb_vpn_12 <= io_tlb12_vpn_i;
    tlb_vpn_13 <= io_tlb13_vpn_i;
    tlb_vpn_14 <= io_tlb14_vpn_i;
    tlb_vpn_15 <= io_tlb15_vpn_i;
    tlb_pte_0 <= io_tlb0_pte_i;
    tlb_pte_1 <= io_tlb1_pte_i;
    tlb_pte_2 <= io_tlb2_pte_i;
    tlb_pte_3 <= io_tlb3_pte_i;
    tlb_pte_4 <= io_tlb4_pte_i;
    tlb_pte_5 <= io_tlb5_pte_i;
    tlb_pte_6 <= io_tlb6_pte_i;
    tlb_pte_7 <= io_tlb7_pte_i;
    tlb_pte_8 <= io_tlb8_pte_i;
    tlb_pte_9 <= io_tlb9_pte_i;
    tlb_pte_10 <= io_tlb10_pte_i;
    tlb_pte_11 <= io_tlb11_pte_i;
    tlb_pte_12 <= io_tlb12_pte_i;
    tlb_pte_13 <= io_tlb13_pte_i;
    tlb_pte_14 <= io_tlb14_pte_i;
    tlb_pte_15 <= io_tlb15_pte_i;
    tlb_mask_0 <= io_tlb0_mask_i;
    tlb_mask_1 <= io_tlb1_mask_i;
    tlb_mask_2 <= io_tlb2_mask_i;
    tlb_mask_3 <= io_tlb3_mask_i;
    tlb_mask_4 <= io_tlb4_mask_i;
    tlb_mask_5 <= io_tlb5_mask_i;
    tlb_mask_6 <= io_tlb6_mask_i;
    tlb_mask_7 <= io_tlb7_mask_i;
    tlb_mask_8 <= io_tlb8_mask_i;
    tlb_mask_9 <= io_tlb9_mask_i;
    tlb_mask_10 <= io_tlb10_mask_i;
    tlb_mask_11 <= io_tlb11_mask_i;
    tlb_mask_12 <= io_tlb12_mask_i;
    tlb_mask_13 <= io_tlb13_mask_i;
    tlb_mask_14 <= io_tlb14_mask_i;
    tlb_mask_15 <= io_tlb15_mask_i;
    phy_addr_0 <= _T_30 | _GEN_287;
    phy_addr_1 <= _T_64 | _GEN_289;
    phy_addr_2 <= _T_98 | _GEN_291;
    phy_addr_3 <= _T_132 | _GEN_293;
    phy_addr_4 <= _T_166 | _GEN_295;
    phy_addr_5 <= _T_200 | _GEN_297;
    phy_addr_6 <= _T_234 | _GEN_299;
    phy_addr_7 <= _T_268 | _GEN_301;
    phy_addr_8 <= _T_302 | _GEN_303;
    phy_addr_9 <= _T_336 | _GEN_305;
    phy_addr_10 <= _T_370 | _GEN_307;
    phy_addr_11 <= _T_404 | _GEN_309;
    phy_addr_12 <= _T_438 | _GEN_311;
    phy_addr_13 <= _T_472 | _GEN_313;
    phy_addr_14 <= _T_506 | _GEN_315;
    phy_addr_15 <= _T_540 | _GEN_317;
  end
endmodule
module CSR(
  input         io_clk,
  input         io_rst_n,
  input         io_we_i,
  input  [11:0] io_waddr_i,
  input  [31:0] io_data_i,
  input         io_re_i,
  input         io_will_write_in_mem_i,
  input  [11:0] io_raddr_i,
  output [31:0] io_data_o,
  output        io_protect_o,
  input         io_inst_ce_i,
  input  [31:0] io_inst_vir_addr_i,
  output [33:0] io_inst_phy_addr_o,
  output        io_inst_tlb_exception_o,
  input         io_data_ce_i,
  input         io_data_we_i,
  input  [31:0] io_data_vir_addr_i,
  output [33:0] io_data_phy_addr_o,
  output        io_data_tlb_exception_o,
  input  [31:0] io_excepttype_i,
  input         io_timer_int_i,
  input         io_external_int_i,
  input         io_software_int_i,
  input  [31:0] io_current_inst_addr_i,
  input  [31:0] io_current_data_addr_i,
  input         io_not_stall_i,
  input         io_is_in_delayslot_i,
  output        io_flushreq,
  output [31:0] io_exception_new_pc_o,
  output [1:0]  io_prv_o
);
  reg [31:0] mtlbvpn [0:15]; // @[CSR.scala 121:26]
  reg [31:0] _RAND_0;
  wire [31:0] mtlbvpn__T_480_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_480_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_483_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_483_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_486_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_486_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_489_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_489_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_492_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_492_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_495_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_495_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_498_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_498_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_501_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_501_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_504_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_504_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_507_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_507_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_510_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_510_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_513_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_513_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_516_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_516_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_519_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_519_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_522_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_522_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_525_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_525_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_528_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_528_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_531_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_531_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_534_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_534_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_537_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_537_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_540_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_540_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_543_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_543_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_546_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_546_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_549_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_549_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_552_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_552_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_555_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_555_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_558_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_558_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_561_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_561_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_564_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_564_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_567_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_567_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_570_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_570_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_573_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_573_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_753_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_753_addr; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_192_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_192_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_192_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_192_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_196_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_196_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_196_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_196_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_200_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_200_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_200_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_200_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_204_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_204_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_204_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_204_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_208_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_208_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_208_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_208_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_212_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_212_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_212_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_212_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_216_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_216_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_216_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_216_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_220_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_220_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_220_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_220_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_224_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_224_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_224_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_224_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_228_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_228_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_228_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_228_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_232_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_232_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_232_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_232_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_236_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_236_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_236_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_236_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_240_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_240_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_240_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_240_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_244_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_244_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_244_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_244_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_248_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_248_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_248_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_248_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_252_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_252_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_252_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_252_en; // @[CSR.scala 121:26]
  wire [31:0] mtlbvpn__T_469_data; // @[CSR.scala 121:26]
  wire [3:0] mtlbvpn__T_469_addr; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_469_mask; // @[CSR.scala 121:26]
  wire  mtlbvpn__T_469_en; // @[CSR.scala 121:26]
  reg [31:0] mtlbmask [0:15]; // @[CSR.scala 122:26]
  reg [31:0] _RAND_1;
  wire [31:0] mtlbmask__T_482_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_482_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_485_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_485_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_488_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_488_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_491_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_491_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_494_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_494_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_497_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_497_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_500_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_500_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_503_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_503_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_506_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_506_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_509_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_509_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_512_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_512_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_515_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_515_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_518_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_518_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_521_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_521_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_524_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_524_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_527_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_527_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_530_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_530_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_533_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_533_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_536_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_536_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_539_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_539_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_542_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_542_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_545_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_545_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_548_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_548_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_551_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_551_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_554_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_554_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_557_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_557_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_560_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_560_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_563_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_563_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_566_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_566_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_569_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_569_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_572_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_572_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_575_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_575_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_755_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_755_addr; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_193_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_193_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_193_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_193_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_197_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_197_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_197_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_197_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_201_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_201_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_201_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_201_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_205_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_205_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_205_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_205_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_209_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_209_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_209_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_209_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_213_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_213_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_213_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_213_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_217_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_217_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_217_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_217_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_221_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_221_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_221_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_221_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_225_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_225_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_225_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_225_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_229_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_229_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_229_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_229_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_233_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_233_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_233_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_233_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_237_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_237_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_237_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_237_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_241_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_241_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_241_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_241_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_245_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_245_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_245_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_245_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_249_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_249_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_249_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_249_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_253_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_253_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_253_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_253_en; // @[CSR.scala 122:26]
  wire [31:0] mtlbmask__T_471_data; // @[CSR.scala 122:26]
  wire [3:0] mtlbmask__T_471_addr; // @[CSR.scala 122:26]
  wire  mtlbmask__T_471_mask; // @[CSR.scala 122:26]
  wire  mtlbmask__T_471_en; // @[CSR.scala 122:26]
  reg [31:0] mtlbpte [0:15]; // @[CSR.scala 123:26]
  reg [31:0] _RAND_2;
  wire [31:0] mtlbpte__T_481_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_481_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_484_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_484_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_487_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_487_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_490_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_490_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_493_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_493_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_496_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_496_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_499_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_499_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_502_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_502_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_505_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_505_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_508_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_508_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_511_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_511_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_514_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_514_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_517_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_517_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_520_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_520_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_523_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_523_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_526_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_526_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_529_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_529_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_532_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_532_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_535_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_535_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_538_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_538_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_541_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_541_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_544_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_544_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_547_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_547_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_550_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_550_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_553_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_553_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_556_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_556_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_559_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_559_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_562_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_562_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_565_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_565_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_568_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_568_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_571_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_571_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_574_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_574_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_757_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_757_addr; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_194_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_194_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_194_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_194_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_198_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_198_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_198_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_198_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_202_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_202_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_202_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_202_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_206_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_206_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_206_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_206_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_210_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_210_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_210_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_210_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_214_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_214_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_214_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_214_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_218_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_218_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_218_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_218_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_222_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_222_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_222_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_222_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_226_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_226_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_226_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_226_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_230_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_230_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_230_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_230_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_234_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_234_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_234_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_234_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_238_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_238_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_238_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_238_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_242_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_242_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_242_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_242_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_246_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_246_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_246_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_246_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_250_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_250_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_250_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_250_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_254_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_254_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_254_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_254_en; // @[CSR.scala 123:26]
  wire [31:0] mtlbpte__T_473_data; // @[CSR.scala 123:26]
  wire [3:0] mtlbpte__T_473_addr; // @[CSR.scala 123:26]
  wire  mtlbpte__T_473_mask; // @[CSR.scala 123:26]
  wire  mtlbpte__T_473_en; // @[CSR.scala 123:26]
  reg [31:0] mtlbptevaddr [0:15]; // @[CSR.scala 124:26]
  reg [31:0] _RAND_3;
  wire [31:0] mtlbptevaddr__T_759_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_759_addr; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_195_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_195_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_195_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_195_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_199_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_199_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_199_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_199_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_203_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_203_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_203_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_203_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_207_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_207_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_207_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_207_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_211_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_211_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_211_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_211_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_215_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_215_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_215_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_215_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_219_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_219_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_219_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_219_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_223_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_223_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_223_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_223_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_227_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_227_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_227_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_227_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_231_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_231_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_231_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_231_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_235_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_235_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_235_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_235_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_239_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_239_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_239_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_239_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_243_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_243_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_243_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_243_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_247_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_247_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_247_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_247_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_251_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_251_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_251_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_251_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_255_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_255_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_255_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_255_en; // @[CSR.scala 124:26]
  wire [31:0] mtlbptevaddr__T_475_data; // @[CSR.scala 124:26]
  wire [3:0] mtlbptevaddr__T_475_addr; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_475_mask; // @[CSR.scala 124:26]
  wire  mtlbptevaddr__T_475_en; // @[CSR.scala 124:26]
  wire  mmu_conv0_clock; // @[CSR.scala 763:25]
  wire  mmu_conv0_io_rst_n; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb0_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb0_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb0_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb1_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb1_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb1_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb2_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb2_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb2_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb3_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb3_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb3_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb4_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb4_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb4_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb5_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb5_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb5_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb6_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb6_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb6_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb7_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb7_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb7_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb8_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb8_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb8_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb9_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb9_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb9_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb10_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb10_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb10_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb11_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb11_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb11_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb12_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb12_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb12_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb13_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb13_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb13_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb14_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb14_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb14_pte_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb15_vpn_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb15_mask_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_tlb15_pte_i; // @[CSR.scala 763:25]
  wire [4:0] mmu_conv0_io_vm_i; // @[CSR.scala 763:25]
  wire [1:0] mmu_conv0_io_prv_i; // @[CSR.scala 763:25]
  wire  mmu_conv0_io_mxr_i; // @[CSR.scala 763:25]
  wire  mmu_conv0_io_ce_i; // @[CSR.scala 763:25]
  wire  mmu_conv0_io_ex_i; // @[CSR.scala 763:25]
  wire  mmu_conv0_io_we_i; // @[CSR.scala 763:25]
  wire [31:0] mmu_conv0_io_vir_addr_i; // @[CSR.scala 763:25]
  wire [33:0] mmu_conv0_io_phy_addr_o; // @[CSR.scala 763:25]
  wire  mmu_conv0_io_tlb_exception_o; // @[CSR.scala 763:25]
  wire  mmu_conv0_io_tlb_update_o; // @[CSR.scala 763:25]
  wire [3:0] mmu_conv0_io_hit_index_o; // @[CSR.scala 763:25]
  wire  mmu_conv1_clock; // @[CSR.scala 799:25]
  wire  mmu_conv1_io_rst_n; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb0_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb0_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb0_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb1_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb1_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb1_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb2_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb2_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb2_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb3_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb3_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb3_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb4_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb4_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb4_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb5_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb5_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb5_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb6_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb6_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb6_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb7_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb7_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb7_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb8_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb8_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb8_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb9_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb9_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb9_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb10_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb10_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb10_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb11_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb11_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb11_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb12_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb12_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb12_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb13_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb13_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb13_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb14_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb14_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb14_pte_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb15_vpn_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb15_mask_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_tlb15_pte_i; // @[CSR.scala 799:25]
  wire [4:0] mmu_conv1_io_vm_i; // @[CSR.scala 799:25]
  wire [1:0] mmu_conv1_io_prv_i; // @[CSR.scala 799:25]
  wire  mmu_conv1_io_mxr_i; // @[CSR.scala 799:25]
  wire  mmu_conv1_io_ce_i; // @[CSR.scala 799:25]
  wire  mmu_conv1_io_ex_i; // @[CSR.scala 799:25]
  wire  mmu_conv1_io_we_i; // @[CSR.scala 799:25]
  wire [31:0] mmu_conv1_io_vir_addr_i; // @[CSR.scala 799:25]
  wire [33:0] mmu_conv1_io_phy_addr_o; // @[CSR.scala 799:25]
  wire  mmu_conv1_io_tlb_exception_o; // @[CSR.scala 799:25]
  wire  mmu_conv1_io_tlb_update_o; // @[CSR.scala 799:25]
  wire [3:0] mmu_conv1_io_hit_index_o; // @[CSR.scala 799:25]
  reg [4:0] mstatus_vm; // @[CSR.scala 72:26]
  reg [31:0] _RAND_4;
  reg  mstatus_mxr; // @[CSR.scala 73:26]
  reg [31:0] _RAND_5;
  reg  mstatus_mprv; // @[CSR.scala 74:26]
  reg [31:0] _RAND_6;
  reg [1:0] mstatus_fs; // @[CSR.scala 75:26]
  reg [31:0] _RAND_7;
  wire  _T_1; // @[CSR.scala 76:53]
  reg  mstatus_sd; // @[CSR.scala 76:30]
  reg [31:0] _RAND_8;
  reg [1:0] mstatus_mpp; // @[CSR.scala 77:26]
  reg [31:0] _RAND_9;
  reg  mstatus_spp; // @[CSR.scala 78:26]
  reg [31:0] _RAND_10;
  reg  mstatus_mpie; // @[CSR.scala 79:26]
  reg [31:0] _RAND_11;
  reg  mstatus_spie; // @[CSR.scala 80:26]
  reg [31:0] _RAND_12;
  reg  mstatus_mie; // @[CSR.scala 81:26]
  reg [31:0] _RAND_13;
  reg  mstatus_sie; // @[CSR.scala 82:26]
  reg [31:0] _RAND_14;
  reg  mip_mtip; // @[CSR.scala 85:27]
  reg [31:0] _RAND_15;
  reg  mip_stip; // @[CSR.scala 86:23]
  reg [31:0] _RAND_16;
  reg  mie_mtie; // @[CSR.scala 87:23]
  reg [31:0] _RAND_17;
  reg  mie_stie; // @[CSR.scala 88:23]
  reg [31:0] _RAND_18;
  reg  mip_msip; // @[CSR.scala 89:27]
  reg [31:0] _RAND_19;
  reg  mip_ssip; // @[CSR.scala 90:23]
  reg [31:0] _RAND_20;
  reg  mie_msie; // @[CSR.scala 91:23]
  reg [31:0] _RAND_21;
  reg  mie_ssie; // @[CSR.scala 92:23]
  reg [31:0] _RAND_22;
  reg  mip_meip; // @[CSR.scala 93:27]
  reg [31:0] _RAND_23;
  reg  mie_meie; // @[CSR.scala 94:23]
  reg [31:0] _RAND_24;
  reg  mucounteren_tm; // @[CSR.scala 96:29]
  reg [31:0] _RAND_25;
  reg  mscounteren_tm; // @[CSR.scala 97:29]
  reg [31:0] _RAND_26;
  reg [31:0] mscratch; // @[CSR.scala 99:24]
  reg [31:0] _RAND_27;
  reg [29:0] mepc_addr; // @[CSR.scala 100:24]
  reg [31:0] _RAND_28;
  reg [29:0] mtvec_addr; // @[CSR.scala 102:24]
  reg [31:0] _RAND_29;
  reg [11:0] medeleg; // @[CSR.scala 103:24]
  reg [31:0] _RAND_30;
  reg [11:0] mideleg; // @[CSR.scala 104:24]
  reg [31:0] _RAND_31;
  reg  mcause_intr; // @[CSR.scala 106:24]
  reg [31:0] _RAND_32;
  reg [3:0] mcause_code; // @[CSR.scala 107:24]
  reg [31:0] _RAND_33;
  reg [31:0] mbadaddr; // @[CSR.scala 108:24]
  reg [31:0] _RAND_34;
  reg [29:0] stvec_addr; // @[CSR.scala 110:24]
  reg [31:0] _RAND_35;
  reg [31:0] sscratch; // @[CSR.scala 111:24]
  reg [31:0] _RAND_36;
  reg [29:0] sepc_addr; // @[CSR.scala 112:24]
  reg [31:0] _RAND_37;
  reg  scause_intr; // @[CSR.scala 113:24]
  reg [31:0] _RAND_38;
  reg [3:0] scause_code; // @[CSR.scala 114:24]
  reg [31:0] _RAND_39;
  reg [31:0] sbadaddr; // @[CSR.scala 115:24]
  reg [31:0] _RAND_40;
  reg [21:0] sptbr_ppn; // @[CSR.scala 117:24]
  reg [31:0] _RAND_41;
  reg [3:0] mtlbindex; // @[CSR.scala 119:30]
  reg [31:0] _RAND_42;
  reg  mtlbindex_update; // @[CSR.scala 120:30]
  reg [31:0] _RAND_43;
  reg [3:0] inst_tlb_index; // @[CSR.scala 126:31]
  reg [31:0] _RAND_44;
  reg  inst_tlb_update; // @[CSR.scala 127:31]
  reg [31:0] _RAND_45;
  reg  inst_tlb_exception; // @[CSR.scala 128:31]
  reg [31:0] _RAND_46;
  reg [3:0] data_tlb_index; // @[CSR.scala 129:31]
  reg [31:0] _RAND_47;
  reg  data_tlb_update; // @[CSR.scala 130:31]
  reg [31:0] _RAND_48;
  reg  data_tlb_exception; // @[CSR.scala 131:31]
  reg [31:0] _RAND_49;
  wire  _T_3; // @[CSR.scala 135:19]
  wire  _T_4; // @[CSR.scala 135:47]
  wire  _T_6; // @[CSR.scala 135:63]
  wire  _T_7; // @[CSR.scala 135:34]
  wire  m_intr_globally_enabled; // @[CSR.scala 135:5]
  wire  _T_9; // @[CSR.scala 140:19]
  wire  _T_10; // @[CSR.scala 140:47]
  wire  _T_12; // @[CSR.scala 140:63]
  wire  _T_13; // @[CSR.scala 140:34]
  wire  s_intr_globally_enabled; // @[CSR.scala 140:5]
  wire  _T_14; // @[CSR.scala 144:31]
  wire  _T_15; // @[CSR.scala 144:42]
  wire  m_mtime_intr; // @[CSR.scala 144:75]
  wire  _T_18; // @[CSR.scala 145:31]
  wire  _T_19; // @[CSR.scala 145:42]
  wire  m_msoft_intr; // @[CSR.scala 145:75]
  wire  _T_22; // @[CSR.scala 146:31]
  wire  _T_23; // @[CSR.scala 146:42]
  wire  m_mextr_intr; // @[CSR.scala 146:75]
  wire  _T_26; // @[CSR.scala 147:31]
  wire  _T_27; // @[CSR.scala 147:42]
  wire  m_stime_intr; // @[CSR.scala 147:75]
  wire  _T_30; // @[CSR.scala 148:31]
  wire  _T_31; // @[CSR.scala 148:42]
  wire  m_ssoft_intr; // @[CSR.scala 148:75]
  wire  _T_34; // @[CSR.scala 150:29]
  wire  _T_35; // @[CSR.scala 150:44]
  wire  _T_36; // @[CSR.scala 150:59]
  wire  m_intr; // @[CSR.scala 150:74]
  wire  _T_38; // @[CSR.scala 152:42]
  wire  s_mtime_intr; // @[CSR.scala 152:75]
  wire  _T_41; // @[CSR.scala 153:42]
  wire  s_msoft_intr; // @[CSR.scala 153:75]
  wire  _T_44; // @[CSR.scala 154:42]
  wire  s_mextr_intr; // @[CSR.scala 154:75]
  wire  _T_47; // @[CSR.scala 155:42]
  wire  s_stime_intr; // @[CSR.scala 155:75]
  wire  _T_50; // @[CSR.scala 156:42]
  wire  s_ssoft_intr; // @[CSR.scala 156:75]
  wire  _T_52; // @[CSR.scala 158:29]
  wire  _T_53; // @[CSR.scala 158:44]
  wire  _T_54; // @[CSR.scala 158:59]
  wire  s_intr; // @[CSR.scala 158:74]
  wire  _T_57; // @[CSR.scala 160:60]
  wire  m_inst_misaligned_trap; // @[CSR.scala 160:110]
  wire [31:0] _T_60; // @[CSR.scala 162:77]
  wire  _T_62; // @[CSR.scala 162:60]
  wire  m_inst_access_fault_trap; // @[CSR.scala 162:110]
  wire [31:0] _T_65; // @[CSR.scala 164:77]
  wire  _T_67; // @[CSR.scala 164:60]
  wire  m_inst_illegal_trap; // @[CSR.scala 164:110]
  wire [31:0] _T_70; // @[CSR.scala 166:77]
  wire  _T_72; // @[CSR.scala 166:60]
  wire  m_break_trap; // @[CSR.scala 166:110]
  wire [31:0] _T_75; // @[CSR.scala 168:77]
  wire  _T_77; // @[CSR.scala 168:60]
  wire  m_load_misaligned_trap; // @[CSR.scala 168:110]
  wire [31:0] _T_80; // @[CSR.scala 170:77]
  wire  _T_82; // @[CSR.scala 170:60]
  wire  m_load_access_fault_trap; // @[CSR.scala 170:110]
  wire [31:0] _T_85; // @[CSR.scala 172:77]
  wire  _T_87; // @[CSR.scala 172:60]
  wire  m_store_misaligned_trap; // @[CSR.scala 172:110]
  wire [31:0] _T_90; // @[CSR.scala 174:77]
  wire  _T_92; // @[CSR.scala 174:60]
  wire  m_store_access_fault_trap; // @[CSR.scala 174:110]
  wire [31:0] _T_95; // @[CSR.scala 176:77]
  wire  _T_97; // @[CSR.scala 176:60]
  wire  m_ecall_from_u_trap; // @[CSR.scala 176:110]
  wire [31:0] _T_100; // @[CSR.scala 178:77]
  wire  _T_102; // @[CSR.scala 178:60]
  wire  m_ecall_from_s_trap; // @[CSR.scala 178:110]
  wire [31:0] _T_105; // @[CSR.scala 180:77]
  wire  m_ecall_from_m_trap; // @[CSR.scala 180:60]
  wire  _T_107; // @[CSR.scala 183:30]
  wire  _T_108; // @[CSR.scala 184:32]
  wire  _T_109; // @[CSR.scala 185:27]
  wire  _T_110; // @[CSR.scala 186:20]
  wire  _T_111; // @[CSR.scala 187:30]
  wire  _T_112; // @[CSR.scala 188:32]
  wire  _T_113; // @[CSR.scala 189:31]
  wire  _T_114; // @[CSR.scala 190:33]
  wire  _T_115; // @[CSR.scala 191:27]
  wire  m_trap; // @[CSR.scala 192:27]
  wire [31:0] _T_116; // @[CSR.scala 195:67]
  wire  eret_from_m_trap; // @[CSR.scala 195:50]
  wire [31:0] _T_118; // @[CSR.scala 196:67]
  wire  eret_from_s_trap; // @[CSR.scala 196:50]
  wire [31:0] _T_120; // @[CSR.scala 197:67]
  wire  fence_i_trap; // @[CSR.scala 197:50]
  wire  s_inst_misaligned_trap; // @[CSR.scala 199:110]
  wire  s_inst_access_fault_trap; // @[CSR.scala 201:110]
  wire  s_inst_illegal_trap; // @[CSR.scala 203:110]
  wire  s_break_trap; // @[CSR.scala 205:110]
  wire  s_load_misaligned_trap; // @[CSR.scala 207:110]
  wire  s_load_access_fault_trap; // @[CSR.scala 209:110]
  wire  s_store_misaligned_trap; // @[CSR.scala 211:110]
  wire  s_store_access_fault_trap; // @[CSR.scala 213:110]
  wire  s_ecall_from_u_trap; // @[CSR.scala 215:110]
  wire  s_ecall_from_s_trap; // @[CSR.scala 217:110]
  wire  _T_162; // @[CSR.scala 220:30]
  wire  _T_163; // @[CSR.scala 221:32]
  wire  _T_164; // @[CSR.scala 222:27]
  wire  _T_165; // @[CSR.scala 223:20]
  wire  _T_166; // @[CSR.scala 224:30]
  wire  _T_167; // @[CSR.scala 225:32]
  wire  _T_168; // @[CSR.scala 226:31]
  wire  _T_169; // @[CSR.scala 227:33]
  wire  s_trap; // @[CSR.scala 228:27]
  reg [1:0] next_prv; // @[CSR.scala 236:21]
  reg [31:0] _RAND_50;
  wire [30:0] _T_172; // @[Cat.scala 29:58]
  wire [30:0] _T_174; // @[Cat.scala 29:58]
  wire [30:0] _T_180; // @[Cat.scala 29:58]
  wire [1:0] _GEN_2048; // @[Conditional.scala 37:30]
  wire  _T_181; // @[Conditional.scala 37:30]
  wire  _T_182; // @[Conditional.scala 37:30]
  wire [30:0] _T_184; // @[Cat.scala 29:58]
  wire  _T_185; // @[Conditional.scala 37:30]
  wire  _T_186; // @[Conditional.scala 37:30]
  wire  _T_187; // @[Conditional.scala 37:30]
  wire [31:0] _T_190; // @[CSR.scala 277:55]
  wire [31:0] _GEN_6; // @[CSR.scala 275:36]
  wire  _GEN_7; // @[CSR.scala 267:40]
  wire [31:0] _GEN_8; // @[CSR.scala 267:40]
  wire  _GEN_10; // @[CSR.scala 260:40]
  wire [31:0] _GEN_11; // @[CSR.scala 260:40]
  wire  _GEN_13; // @[CSR.scala 256:30]
  wire [31:0] _GEN_14; // @[CSR.scala 256:30]
  wire  _GEN_16; // @[CSR.scala 252:30]
  wire [31:0] _GEN_17; // @[CSR.scala 252:30]
  wire  _GEN_19; // @[CSR.scala 248:30]
  wire [31:0] _GEN_20; // @[CSR.scala 248:30]
  wire  _GEN_22; // @[CSR.scala 244:24]
  wire [31:0] _GEN_23; // @[CSR.scala 244:24]
  wire  _GEN_28; // @[CSR.scala 365:37]
  wire [3:0] _GEN_29; // @[CSR.scala 365:37]
  wire  _GEN_30; // @[CSR.scala 362:37]
  wire [3:0] _GEN_31; // @[CSR.scala 362:37]
  wire  _GEN_32; // @[CSR.scala 359:37]
  wire [3:0] _GEN_33; // @[CSR.scala 359:37]
  wire  _GEN_34; // @[CSR.scala 356:37]
  wire [3:0] _GEN_35; // @[CSR.scala 356:37]
  wire  _GEN_36; // @[CSR.scala 353:31]
  wire [3:0] _GEN_37; // @[CSR.scala 353:31]
  wire  _T_264; // @[Conditional.scala 37:30]
  wire  _T_265; // @[Conditional.scala 37:30]
  wire  _T_266; // @[Conditional.scala 37:30]
  wire  _GEN_44; // @[CSR.scala 399:37]
  wire [3:0] _GEN_45; // @[CSR.scala 399:37]
  wire  _GEN_46; // @[CSR.scala 396:37]
  wire [3:0] _GEN_47; // @[CSR.scala 396:37]
  wire  _GEN_48; // @[CSR.scala 393:37]
  wire [3:0] _GEN_49; // @[CSR.scala 393:37]
  wire  _GEN_50; // @[CSR.scala 390:37]
  wire [3:0] _GEN_51; // @[CSR.scala 390:37]
  wire  _GEN_52; // @[CSR.scala 387:31]
  wire [3:0] _GEN_53; // @[CSR.scala 387:31]
  wire [1:0] _GEN_56; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_57; // @[Conditional.scala 40:58]
  wire [3:0] _GEN_59; // @[CSR.scala 455:44]
  wire [3:0] _GEN_61; // @[CSR.scala 452:44]
  wire [3:0] _GEN_63; // @[CSR.scala 449:44]
  wire [3:0] _GEN_65; // @[CSR.scala 445:50]
  wire [3:0] _GEN_68; // @[CSR.scala 441:48]
  wire [3:0] _GEN_71; // @[CSR.scala 437:49]
  wire [3:0] _GEN_74; // @[CSR.scala 433:47]
  wire [3:0] _GEN_77; // @[CSR.scala 430:37]
  wire [3:0] _GEN_80; // @[CSR.scala 427:44]
  wire [3:0] _GEN_83; // @[CSR.scala 423:49]
  wire [3:0] _GEN_86; // @[CSR.scala 419:41]
  wire [3:0] _GEN_95; // @[CSR.scala 510:44]
  wire [3:0] _GEN_97; // @[CSR.scala 507:44]
  wire [3:0] _GEN_99; // @[CSR.scala 503:50]
  wire [3:0] _GEN_102; // @[CSR.scala 499:48]
  wire [3:0] _GEN_105; // @[CSR.scala 495:49]
  wire [3:0] _GEN_108; // @[CSR.scala 491:47]
  wire [3:0] _GEN_111; // @[CSR.scala 488:37]
  wire [3:0] _GEN_114; // @[CSR.scala 485:44]
  wire [3:0] _GEN_117; // @[CSR.scala 481:49]
  wire [3:0] _GEN_120; // @[CSR.scala 477:41]
  wire  _GEN_127; // @[Conditional.scala 39:67]
  wire  _GEN_128; // @[Conditional.scala 39:67]
  wire  _GEN_129; // @[Conditional.scala 40:58]
  wire  _GEN_130; // @[Conditional.scala 40:58]
  wire  _GEN_133; // @[Conditional.scala 39:67]
  wire  _GEN_136; // @[Conditional.scala 39:67]
  wire  _GEN_138; // @[Conditional.scala 40:58]
  wire  _T_325; // @[Conditional.scala 37:30]
  wire  _T_327; // @[Conditional.scala 37:30]
  wire  _T_328; // @[Conditional.scala 37:30]
  wire  _T_329; // @[Conditional.scala 37:55]
  wire  _T_335; // @[Conditional.scala 37:30]
  wire  _T_336; // @[Conditional.scala 37:30]
  wire  _T_337; // @[Conditional.scala 37:30]
  wire  _T_338; // @[Conditional.scala 37:55]
  wire  _T_339; // @[Conditional.scala 37:55]
  wire [1:0] _T_342; // @[Cat.scala 29:58]
  wire  _T_343; // @[Conditional.scala 37:30]
  wire  _T_344; // @[Conditional.scala 37:30]
  wire  _T_345; // @[Conditional.scala 37:55]
  wire  _GEN_143; // @[Conditional.scala 40:58]
  wire  _T_351; // @[Conditional.scala 37:30]
  wire  _T_354; // @[Conditional.scala 37:30]
  wire  _T_360; // @[Conditional.scala 37:30]
  wire  _T_362; // @[Conditional.scala 37:30]
  wire  _T_364; // @[Conditional.scala 37:30]
  wire  _T_365; // @[Conditional.scala 37:30]
  wire  _T_367; // @[Conditional.scala 37:30]
  wire  _T_369; // @[Conditional.scala 37:30]
  wire  _T_371; // @[Conditional.scala 37:30]
  wire  _T_373; // @[Conditional.scala 37:30]
  wire [4:0] _T_376; // @[Cat.scala 29:58]
  wire  _T_377; // @[Conditional.scala 37:30]
  wire  _T_378; // @[Conditional.scala 37:30]
  wire  _T_379; // @[Conditional.scala 37:30]
  wire  _T_380; // @[Conditional.scala 37:30]
  wire  _T_381; // @[Conditional.scala 37:30]
  wire  _T_382; // @[Conditional.scala 37:30]
  wire  _T_383; // @[Conditional.scala 37:30]
  wire  _T_384; // @[Conditional.scala 37:30]
  wire  _T_385; // @[Conditional.scala 37:30]
  wire  _T_386; // @[Conditional.scala 37:30]
  wire  _T_387; // @[Conditional.scala 37:30]
  wire  _T_388; // @[Conditional.scala 37:30]
  wire  _T_389; // @[Conditional.scala 37:30]
  wire  _T_390; // @[Conditional.scala 37:30]
  wire  _T_391; // @[Conditional.scala 37:30]
  wire  _T_392; // @[Conditional.scala 37:30]
  wire  _T_393; // @[Conditional.scala 37:30]
  wire  _T_394; // @[Conditional.scala 37:55]
  wire  _T_395; // @[Conditional.scala 37:55]
  wire  _T_396; // @[Conditional.scala 37:55]
  wire  _T_397; // @[Conditional.scala 37:55]
  wire  _T_398; // @[Conditional.scala 37:55]
  wire  _T_399; // @[Conditional.scala 37:55]
  wire  _T_400; // @[Conditional.scala 37:55]
  wire  _T_401; // @[Conditional.scala 37:55]
  wire  _T_402; // @[Conditional.scala 37:55]
  wire  _T_403; // @[Conditional.scala 37:55]
  wire  _T_404; // @[Conditional.scala 37:55]
  wire  _T_405; // @[Conditional.scala 37:55]
  wire  _T_406; // @[Conditional.scala 37:55]
  wire  _T_407; // @[Conditional.scala 37:55]
  wire  _T_408; // @[Conditional.scala 37:55]
  wire  _T_409; // @[Conditional.scala 37:55]
  wire [3:0] _GEN_145; // @[Conditional.scala 40:58]
  wire  _T_412; // @[Conditional.scala 37:30]
  wire  _T_413; // @[Conditional.scala 37:30]
  wire  _T_423; // @[Conditional.scala 37:30]
  wire  _T_425; // @[Conditional.scala 37:30]
  wire  _T_428; // @[Conditional.scala 37:30]
  wire  _T_431; // @[Conditional.scala 37:30]
  wire  _T_432; // @[Conditional.scala 37:30]
  wire  _T_434; // @[Conditional.scala 37:30]
  wire  _T_459; // @[Conditional.scala 37:55]
  wire  _T_460; // @[Conditional.scala 37:55]
  wire [3:0] _GEN_148; // @[Conditional.scala 40:58]
  wire  _T_463; // @[Conditional.scala 37:30]
  wire  _T_464; // @[Conditional.scala 37:30]
  wire  _T_466; // @[Conditional.scala 37:30]
  wire  _T_468; // @[Conditional.scala 37:30]
  wire  _T_470; // @[Conditional.scala 37:30]
  wire  _T_472; // @[Conditional.scala 37:30]
  wire  _T_474; // @[Conditional.scala 37:30]
  wire  _GEN_161; // @[Conditional.scala 39:67]
  wire  _GEN_171; // @[Conditional.scala 39:67]
  wire  _GEN_176; // @[Conditional.scala 39:67]
  wire  _GEN_186; // @[Conditional.scala 39:67]
  wire  _GEN_191; // @[Conditional.scala 39:67]
  wire  _GEN_196; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_199; // @[Conditional.scala 39:67]
  wire  _GEN_200; // @[Conditional.scala 39:67]
  wire  _GEN_203; // @[Conditional.scala 39:67]
  wire  _GEN_208; // @[Conditional.scala 39:67]
  wire  _GEN_213; // @[Conditional.scala 39:67]
  wire  _GEN_218; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_221; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_222; // @[Conditional.scala 39:67]
  wire  _GEN_223; // @[Conditional.scala 39:67]
  wire  _GEN_226; // @[Conditional.scala 39:67]
  wire  _GEN_231; // @[Conditional.scala 39:67]
  wire  _GEN_236; // @[Conditional.scala 39:67]
  wire  _GEN_241; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_245; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_246; // @[Conditional.scala 39:67]
  wire  _GEN_247; // @[Conditional.scala 39:67]
  wire  _GEN_250; // @[Conditional.scala 39:67]
  wire  _GEN_255; // @[Conditional.scala 39:67]
  wire  _GEN_260; // @[Conditional.scala 39:67]
  wire  _GEN_265; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_269; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_271; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_272; // @[Conditional.scala 39:67]
  wire  _GEN_273; // @[Conditional.scala 39:67]
  wire  _GEN_276; // @[Conditional.scala 39:67]
  wire  _GEN_281; // @[Conditional.scala 39:67]
  wire  _GEN_286; // @[Conditional.scala 39:67]
  wire  _GEN_291; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_294; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_296; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_298; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_299; // @[Conditional.scala 39:67]
  wire  _GEN_300; // @[Conditional.scala 39:67]
  wire  _GEN_303; // @[Conditional.scala 39:67]
  wire  _GEN_308; // @[Conditional.scala 39:67]
  wire  _GEN_313; // @[Conditional.scala 39:67]
  wire  _GEN_318; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_322; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_324; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_326; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_327; // @[Conditional.scala 39:67]
  wire  _GEN_328; // @[Conditional.scala 39:67]
  wire  _GEN_331; // @[Conditional.scala 39:67]
  wire  _GEN_336; // @[Conditional.scala 39:67]
  wire  _GEN_341; // @[Conditional.scala 39:67]
  wire  _GEN_346; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_352; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_354; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_356; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_357; // @[Conditional.scala 39:67]
  wire  _GEN_358; // @[Conditional.scala 39:67]
  wire  _GEN_361; // @[Conditional.scala 39:67]
  wire  _GEN_366; // @[Conditional.scala 39:67]
  wire  _GEN_371; // @[Conditional.scala 39:67]
  wire  _GEN_376; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_384; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_386; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_388; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_389; // @[Conditional.scala 39:67]
  wire  _GEN_390; // @[Conditional.scala 39:67]
  wire  _GEN_393; // @[Conditional.scala 39:67]
  wire  _GEN_398; // @[Conditional.scala 39:67]
  wire  _GEN_403; // @[Conditional.scala 39:67]
  wire  _GEN_408; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_411; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_417; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_419; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_421; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_422; // @[Conditional.scala 39:67]
  wire  _GEN_423; // @[Conditional.scala 39:67]
  wire  _GEN_426; // @[Conditional.scala 39:67]
  wire  _GEN_431; // @[Conditional.scala 39:67]
  wire  _GEN_436; // @[Conditional.scala 39:67]
  wire  _GEN_441; // @[Conditional.scala 39:67]
  wire  _GEN_445; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_448; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_454; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_456; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_458; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_459; // @[Conditional.scala 39:67]
  wire  _GEN_460; // @[Conditional.scala 39:67]
  wire  _GEN_463; // @[Conditional.scala 39:67]
  wire  _GEN_468; // @[Conditional.scala 39:67]
  wire  _GEN_473; // @[Conditional.scala 39:67]
  wire  _GEN_478; // @[Conditional.scala 39:67]
  wire  _GEN_483; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_486; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_492; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_494; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_496; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_497; // @[Conditional.scala 39:67]
  wire  _GEN_498; // @[Conditional.scala 39:67]
  wire  _GEN_501; // @[Conditional.scala 39:67]
  wire  _GEN_506; // @[Conditional.scala 39:67]
  wire  _GEN_511; // @[Conditional.scala 39:67]
  wire  _GEN_516; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_520; // @[Conditional.scala 39:67]
  wire  _GEN_523; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_526; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_532; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_534; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_536; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_537; // @[Conditional.scala 39:67]
  wire  _GEN_538; // @[Conditional.scala 39:67]
  wire  _GEN_541; // @[Conditional.scala 39:67]
  wire  _GEN_546; // @[Conditional.scala 39:67]
  wire  _GEN_551; // @[Conditional.scala 39:67]
  wire  _GEN_556; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_559; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_561; // @[Conditional.scala 39:67]
  wire  _GEN_564; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_567; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_573; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_575; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_577; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_578; // @[Conditional.scala 39:67]
  wire  _GEN_579; // @[Conditional.scala 39:67]
  wire  _GEN_582; // @[Conditional.scala 39:67]
  wire  _GEN_587; // @[Conditional.scala 39:67]
  wire  _GEN_592; // @[Conditional.scala 39:67]
  wire  _GEN_597; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_600; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_601; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_603; // @[Conditional.scala 39:67]
  wire  _GEN_606; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_609; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_615; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_617; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_619; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_620; // @[Conditional.scala 39:67]
  wire  _GEN_621; // @[Conditional.scala 39:67]
  wire  _GEN_624; // @[Conditional.scala 39:67]
  wire  _GEN_629; // @[Conditional.scala 39:67]
  wire  _GEN_634; // @[Conditional.scala 39:67]
  wire  _GEN_639; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_642; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_643; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_644; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_646; // @[Conditional.scala 39:67]
  wire  _GEN_649; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_652; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_658; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_660; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_662; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_663; // @[Conditional.scala 39:67]
  wire  _GEN_664; // @[Conditional.scala 39:67]
  wire  _GEN_667; // @[Conditional.scala 39:67]
  wire  _GEN_672; // @[Conditional.scala 39:67]
  wire  _GEN_677; // @[Conditional.scala 39:67]
  wire  _GEN_682; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_685; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_686; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_687; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_688; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_690; // @[Conditional.scala 39:67]
  wire  _GEN_693; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_696; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_702; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_704; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_706; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_707; // @[Conditional.scala 39:67]
  wire  _GEN_708; // @[Conditional.scala 39:67]
  wire  _GEN_711; // @[Conditional.scala 39:67]
  wire  _GEN_716; // @[Conditional.scala 39:67]
  wire  _GEN_721; // @[Conditional.scala 39:67]
  wire  _GEN_726; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_730; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_731; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_732; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_733; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_735; // @[Conditional.scala 39:67]
  wire  _GEN_738; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_741; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_747; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_749; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_751; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_752; // @[Conditional.scala 39:67]
  wire  _GEN_753; // @[Conditional.scala 39:67]
  wire  _GEN_756; // @[Conditional.scala 39:67]
  wire  _GEN_761; // @[Conditional.scala 39:67]
  wire  _GEN_766; // @[Conditional.scala 39:67]
  wire  _GEN_771; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_776; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_777; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_778; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_779; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_781; // @[Conditional.scala 39:67]
  wire  _GEN_784; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_787; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_793; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_795; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_797; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_798; // @[Conditional.scala 39:67]
  wire  _GEN_799; // @[Conditional.scala 39:67]
  wire  _GEN_802; // @[Conditional.scala 39:67]
  wire  _GEN_807; // @[Conditional.scala 39:67]
  wire  _GEN_812; // @[Conditional.scala 39:67]
  wire  _GEN_817; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_823; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_824; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_825; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_826; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_828; // @[Conditional.scala 39:67]
  wire  _GEN_831; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_834; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_840; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_842; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_844; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_845; // @[Conditional.scala 39:67]
  wire  _GEN_846; // @[Conditional.scala 39:67]
  wire  _GEN_849; // @[Conditional.scala 39:67]
  wire  _GEN_854; // @[Conditional.scala 39:67]
  wire  _GEN_859; // @[Conditional.scala 39:67]
  wire  _GEN_864; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_875; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_876; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_877; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_878; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_880; // @[Conditional.scala 39:67]
  wire  _GEN_883; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_886; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_890; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_892; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_894; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_895; // @[Conditional.scala 39:67]
  wire  _GEN_896; // @[Conditional.scala 39:67]
  wire  _GEN_899; // @[Conditional.scala 39:67]
  wire  _GEN_904; // @[Conditional.scala 39:67]
  wire  _GEN_909; // @[Conditional.scala 39:67]
  wire  _GEN_914; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_927; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_928; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_929; // @[Conditional.scala 39:67]
  wire [11:0] _GEN_930; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_932; // @[Conditional.scala 39:67]
  wire  _GEN_935; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_938; // @[Conditional.scala 39:67]
  wire [29:0] _GEN_940; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_942; // @[Conditional.scala 39:67]
  wire [21:0] _GEN_944; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_945; // @[Conditional.scala 39:67]
  wire  _GEN_946; // @[Conditional.scala 39:67]
  wire  _GEN_949; // @[Conditional.scala 39:67]
  wire  _GEN_954; // @[Conditional.scala 39:67]
  wire  _GEN_959; // @[Conditional.scala 39:67]
  wire  _GEN_964; // @[Conditional.scala 39:67]
  wire  _GEN_972; // @[Conditional.scala 40:58]
  wire [29:0] _GEN_987; // @[Conditional.scala 40:58]
  wire [29:0] _GEN_988; // @[Conditional.scala 40:58]
  wire [11:0] _GEN_989; // @[Conditional.scala 40:58]
  wire [11:0] _GEN_990; // @[Conditional.scala 40:58]
  wire [3:0] _GEN_992; // @[Conditional.scala 40:58]
  wire [29:0] _GEN_994; // @[Conditional.scala 40:58]
  wire [29:0] _GEN_996; // @[Conditional.scala 40:58]
  wire [3:0] _GEN_998; // @[Conditional.scala 40:58]
  wire [21:0] _GEN_1000; // @[Conditional.scala 40:58]
  wire [3:0] _GEN_1001; // @[Conditional.scala 40:58]
  wire  _GEN_1002; // @[Conditional.scala 40:58]
  wire  _GEN_1005; // @[Conditional.scala 40:58]
  wire  _GEN_1010; // @[Conditional.scala 40:58]
  wire  _GEN_1015; // @[Conditional.scala 40:58]
  wire  _GEN_1020; // @[Conditional.scala 40:58]
  wire  _GEN_1028; // @[CSR.scala 561:34]
  wire [29:0] _GEN_1043; // @[CSR.scala 561:34]
  wire [29:0] _GEN_1044; // @[CSR.scala 561:34]
  wire [11:0] _GEN_1045; // @[CSR.scala 561:34]
  wire [11:0] _GEN_1046; // @[CSR.scala 561:34]
  wire [3:0] _GEN_1048; // @[CSR.scala 561:34]
  wire [29:0] _GEN_1050; // @[CSR.scala 561:34]
  wire [29:0] _GEN_1052; // @[CSR.scala 561:34]
  wire [3:0] _GEN_1054; // @[CSR.scala 561:34]
  wire [21:0] _GEN_1056; // @[CSR.scala 561:34]
  wire [3:0] _GEN_1057; // @[CSR.scala 561:34]
  wire  _GEN_1058; // @[CSR.scala 561:34]
  wire  _GEN_1061; // @[CSR.scala 561:34]
  wire  _GEN_1066; // @[CSR.scala 561:34]
  wire  _GEN_1071; // @[CSR.scala 561:34]
  wire  _GEN_1076; // @[CSR.scala 561:34]
  wire  _GEN_1084; // @[CSR.scala 559:35]
  wire [29:0] _GEN_1099; // @[CSR.scala 559:35]
  wire [29:0] _GEN_1100; // @[CSR.scala 559:35]
  wire [11:0] _GEN_1101; // @[CSR.scala 559:35]
  wire [11:0] _GEN_1102; // @[CSR.scala 559:35]
  wire [3:0] _GEN_1104; // @[CSR.scala 559:35]
  wire [29:0] _GEN_1106; // @[CSR.scala 559:35]
  wire [29:0] _GEN_1108; // @[CSR.scala 559:35]
  wire [3:0] _GEN_1110; // @[CSR.scala 559:35]
  wire [21:0] _GEN_1112; // @[CSR.scala 559:35]
  wire [3:0] _GEN_1113; // @[CSR.scala 559:35]
  wire  _GEN_1114; // @[CSR.scala 559:35]
  wire  _GEN_1117; // @[CSR.scala 559:35]
  wire  _GEN_1122; // @[CSR.scala 559:35]
  wire  _GEN_1127; // @[CSR.scala 559:35]
  wire  _GEN_1132; // @[CSR.scala 559:35]
  wire  _GEN_1142; // @[CSR.scala 540:39]
  wire [29:0] _GEN_1155; // @[CSR.scala 540:39]
  wire [29:0] _GEN_1156; // @[CSR.scala 540:39]
  wire [11:0] _GEN_1157; // @[CSR.scala 540:39]
  wire [11:0] _GEN_1158; // @[CSR.scala 540:39]
  wire [3:0] _GEN_1160; // @[CSR.scala 540:39]
  wire [29:0] _GEN_1162; // @[CSR.scala 540:39]
  wire [29:0] _GEN_1164; // @[CSR.scala 540:39]
  wire [3:0] _GEN_1166; // @[CSR.scala 540:39]
  wire [21:0] _GEN_1168; // @[CSR.scala 540:39]
  wire [3:0] _GEN_1169; // @[CSR.scala 540:39]
  wire  _GEN_1170; // @[CSR.scala 540:39]
  wire  _GEN_1173; // @[CSR.scala 540:39]
  wire  _GEN_1178; // @[CSR.scala 540:39]
  wire  _GEN_1183; // @[CSR.scala 540:39]
  wire  _GEN_1188; // @[CSR.scala 540:39]
  wire  _GEN_1192; // @[CSR.scala 527:39]
  wire [29:0] _GEN_1211; // @[CSR.scala 527:39]
  wire [29:0] _GEN_1212; // @[CSR.scala 527:39]
  wire [11:0] _GEN_1213; // @[CSR.scala 527:39]
  wire [11:0] _GEN_1214; // @[CSR.scala 527:39]
  wire [3:0] _GEN_1216; // @[CSR.scala 527:39]
  wire [29:0] _GEN_1218; // @[CSR.scala 527:39]
  wire [29:0] _GEN_1220; // @[CSR.scala 527:39]
  wire [3:0] _GEN_1222; // @[CSR.scala 527:39]
  wire [21:0] _GEN_1224; // @[CSR.scala 527:39]
  wire [3:0] _GEN_1225; // @[CSR.scala 527:39]
  wire  _GEN_1226; // @[CSR.scala 527:39]
  wire  _GEN_1229; // @[CSR.scala 527:39]
  wire  _GEN_1234; // @[CSR.scala 527:39]
  wire  _GEN_1239; // @[CSR.scala 527:39]
  wire  _GEN_1244; // @[CSR.scala 527:39]
  wire [29:0] _GEN_1247; // @[CSR.scala 474:29]
  wire [3:0] _GEN_1249; // @[CSR.scala 474:29]
  wire [1:0] _GEN_1252; // @[CSR.scala 474:29]
  wire [29:0] _GEN_1271; // @[CSR.scala 474:29]
  wire [29:0] _GEN_1272; // @[CSR.scala 474:29]
  wire [11:0] _GEN_1273; // @[CSR.scala 474:29]
  wire [11:0] _GEN_1274; // @[CSR.scala 474:29]
  wire [29:0] _GEN_1275; // @[CSR.scala 474:29]
  wire [3:0] _GEN_1278; // @[CSR.scala 474:29]
  wire [21:0] _GEN_1280; // @[CSR.scala 474:29]
  wire [3:0] _GEN_1281; // @[CSR.scala 474:29]
  wire  _GEN_1282; // @[CSR.scala 474:29]
  wire  _GEN_1285; // @[CSR.scala 474:29]
  wire  _GEN_1290; // @[CSR.scala 474:29]
  wire  _GEN_1295; // @[CSR.scala 474:29]
  wire  _GEN_1300; // @[CSR.scala 474:29]
  wire [29:0] _GEN_1303; // @[CSR.scala 416:29]
  wire [3:0] _GEN_1305; // @[CSR.scala 416:29]
  wire [29:0] _GEN_1310; // @[CSR.scala 416:29]
  wire [1:0] _GEN_1312; // @[CSR.scala 416:29]
  wire [29:0] _GEN_1328; // @[CSR.scala 416:29]
  wire [11:0] _GEN_1329; // @[CSR.scala 416:29]
  wire [11:0] _GEN_1330; // @[CSR.scala 416:29]
  wire [29:0] _GEN_1331; // @[CSR.scala 416:29]
  wire [3:0] _GEN_1334; // @[CSR.scala 416:29]
  wire [21:0] _GEN_1336; // @[CSR.scala 416:29]
  wire [3:0] _GEN_1337; // @[CSR.scala 416:29]
  wire  _GEN_1338; // @[CSR.scala 416:29]
  wire  _GEN_1341; // @[CSR.scala 416:29]
  wire  _GEN_1346; // @[CSR.scala 416:29]
  wire  _GEN_1351; // @[CSR.scala 416:29]
  wire  _GEN_1356; // @[CSR.scala 416:29]
  wire [29:0] _GEN_1359; // @[CSR.scala 384:29]
  wire [3:0] _GEN_1361; // @[CSR.scala 384:29]
  wire [1:0] _GEN_1363; // @[CSR.scala 384:29]
  wire [29:0] _GEN_1365; // @[CSR.scala 384:29]
  wire [3:0] _GEN_1367; // @[CSR.scala 384:29]
  wire [29:0] _GEN_1386; // @[CSR.scala 384:29]
  wire [11:0] _GEN_1387; // @[CSR.scala 384:29]
  wire [11:0] _GEN_1388; // @[CSR.scala 384:29]
  wire [29:0] _GEN_1389; // @[CSR.scala 384:29]
  wire [21:0] _GEN_1392; // @[CSR.scala 384:29]
  wire [3:0] _GEN_1393; // @[CSR.scala 384:29]
  wire  _GEN_1394; // @[CSR.scala 384:29]
  wire  _GEN_1397; // @[CSR.scala 384:29]
  wire  _GEN_1402; // @[CSR.scala 384:29]
  wire  _GEN_1407; // @[CSR.scala 384:29]
  wire  _GEN_1412; // @[CSR.scala 384:29]
  wire [29:0] _GEN_1415; // @[CSR.scala 350:29]
  wire [3:0] _GEN_1417; // @[CSR.scala 350:29]
  wire [29:0] _GEN_1421; // @[CSR.scala 350:29]
  wire [3:0] _GEN_1423; // @[CSR.scala 350:29]
  wire [1:0] _GEN_1425; // @[CSR.scala 350:29]
  wire [29:0] _GEN_1442; // @[CSR.scala 350:29]
  wire [11:0] _GEN_1443; // @[CSR.scala 350:29]
  wire [11:0] _GEN_1444; // @[CSR.scala 350:29]
  wire [29:0] _GEN_1445; // @[CSR.scala 350:29]
  wire [21:0] _GEN_1448; // @[CSR.scala 350:29]
  wire [3:0] _GEN_1449; // @[CSR.scala 350:29]
  wire  _GEN_1450; // @[CSR.scala 350:29]
  wire  _GEN_1453; // @[CSR.scala 350:29]
  wire  _GEN_1458; // @[CSR.scala 350:29]
  wire  _GEN_1463; // @[CSR.scala 350:29]
  wire  _GEN_1468; // @[CSR.scala 350:29]
  wire [29:0] _GEN_1471; // @[CSR.scala 348:25]
  wire [3:0] _GEN_1473; // @[CSR.scala 348:25]
  wire [29:0] _GEN_1477; // @[CSR.scala 348:25]
  wire [3:0] _GEN_1479; // @[CSR.scala 348:25]
  wire [1:0] _GEN_1481; // @[CSR.scala 348:25]
  wire [29:0] _GEN_1498; // @[CSR.scala 348:25]
  wire [11:0] _GEN_1499; // @[CSR.scala 348:25]
  wire [11:0] _GEN_1500; // @[CSR.scala 348:25]
  wire [29:0] _GEN_1501; // @[CSR.scala 348:25]
  wire [21:0] _GEN_1504; // @[CSR.scala 348:25]
  wire [3:0] _GEN_1505; // @[CSR.scala 348:25]
  wire  _GEN_1506; // @[CSR.scala 348:25]
  wire  _GEN_1509; // @[CSR.scala 348:25]
  wire  _GEN_1514; // @[CSR.scala 348:25]
  wire  _GEN_1519; // @[CSR.scala 348:25]
  wire  _GEN_1524; // @[CSR.scala 348:25]
  wire  _GEN_1527; // @[CSR.scala 754:41]
  wire [3:0] _GEN_1528; // @[CSR.scala 751:38]
  wire  _GEN_1529; // @[CSR.scala 751:38]
  wire  _GEN_1530; // @[CSR.scala 749:41]
  wire [3:0] _GEN_1531; // @[CSR.scala 749:41]
  wire [3:0] _GEN_1532; // @[CSR.scala 746:32]
  wire  _GEN_1533; // @[CSR.scala 746:32]
  wire [1:0] _GEN_1539; // @[CSR.scala 283:32]
  wire [31:0] _GEN_1554; // @[CSR.scala 283:32]
  wire [31:0] _GEN_1555; // @[CSR.scala 283:32]
  wire [31:0] _GEN_1556; // @[CSR.scala 283:32]
  wire [31:0] _GEN_1557; // @[CSR.scala 283:32]
  wire [31:0] _GEN_1559; // @[CSR.scala 283:32]
  wire [31:0] _GEN_1561; // @[CSR.scala 283:32]
  wire [31:0] _GEN_1563; // @[CSR.scala 283:32]
  wire [31:0] _GEN_1565; // @[CSR.scala 283:32]
  wire [31:0] _GEN_1567; // @[CSR.scala 283:32]
  wire [31:0] _GEN_1568; // @[CSR.scala 283:32]
  wire  _T_582; // @[CSR.scala 838:40]
  wire  _T_584; // @[CSR.scala 840:23]
  wire  _T_587; // @[CSR.scala 842:73]
  wire  _T_588; // @[CSR.scala 842:52]
  wire  _T_589; // @[Conditional.scala 37:30]
  wire  _T_590; // @[Conditional.scala 37:30]
  wire  _T_591; // @[Conditional.scala 37:30]
  wire  _T_592; // @[Conditional.scala 37:30]
  wire  _T_593; // @[Conditional.scala 37:30]
  wire  _T_594; // @[Conditional.scala 37:30]
  wire  _T_595; // @[Conditional.scala 37:30]
  wire  _T_596; // @[Conditional.scala 37:30]
  wire  _T_597; // @[Conditional.scala 37:30]
  wire  _T_598; // @[Conditional.scala 37:30]
  wire  _T_599; // @[Conditional.scala 37:30]
  wire  _T_600; // @[Conditional.scala 37:30]
  wire  _T_601; // @[Conditional.scala 37:30]
  wire  _T_602; // @[Conditional.scala 37:30]
  wire  _T_603; // @[Conditional.scala 37:30]
  wire  _T_604; // @[Conditional.scala 37:30]
  wire  _T_605; // @[Conditional.scala 37:30]
  wire  _T_606; // @[Conditional.scala 37:30]
  wire  _T_607; // @[Conditional.scala 37:30]
  wire  _T_608; // @[Conditional.scala 37:30]
  wire  _T_609; // @[Conditional.scala 37:30]
  wire  _T_610; // @[Conditional.scala 37:30]
  wire  _T_611; // @[Conditional.scala 37:30]
  wire  _T_612; // @[Conditional.scala 37:30]
  wire  _T_613; // @[Conditional.scala 37:30]
  wire  _T_614; // @[Conditional.scala 37:30]
  wire  _T_615; // @[Conditional.scala 37:30]
  wire  _T_616; // @[Conditional.scala 37:30]
  wire  _T_617; // @[Conditional.scala 37:30]
  wire  _T_618; // @[Conditional.scala 37:30]
  wire  _T_619; // @[Conditional.scala 37:30]
  wire  _T_620; // @[Conditional.scala 37:55]
  wire  _T_621; // @[Conditional.scala 37:55]
  wire  _T_622; // @[Conditional.scala 37:55]
  wire  _T_623; // @[Conditional.scala 37:55]
  wire  _T_624; // @[Conditional.scala 37:55]
  wire  _T_625; // @[Conditional.scala 37:55]
  wire  _T_626; // @[Conditional.scala 37:55]
  wire  _T_627; // @[Conditional.scala 37:55]
  wire  _T_628; // @[Conditional.scala 37:55]
  wire  _T_629; // @[Conditional.scala 37:55]
  wire  _T_630; // @[Conditional.scala 37:55]
  wire  _T_631; // @[Conditional.scala 37:55]
  wire  _T_632; // @[Conditional.scala 37:55]
  wire  _T_633; // @[Conditional.scala 37:55]
  wire  _T_634; // @[Conditional.scala 37:55]
  wire  _T_635; // @[Conditional.scala 37:55]
  wire  _T_636; // @[Conditional.scala 37:55]
  wire  _T_637; // @[Conditional.scala 37:55]
  wire  _T_638; // @[Conditional.scala 37:55]
  wire  _T_639; // @[Conditional.scala 37:55]
  wire  _T_640; // @[Conditional.scala 37:55]
  wire  _T_641; // @[Conditional.scala 37:55]
  wire  _T_642; // @[Conditional.scala 37:55]
  wire  _T_643; // @[Conditional.scala 37:55]
  wire  _T_644; // @[Conditional.scala 37:55]
  wire  _T_645; // @[Conditional.scala 37:55]
  wire  _T_646; // @[Conditional.scala 37:55]
  wire  _T_647; // @[Conditional.scala 37:55]
  wire  _T_648; // @[Conditional.scala 37:55]
  wire  _T_649; // @[Conditional.scala 37:55]
  wire  _GEN_1611; // @[CSR.scala 842:90]
  wire  _GEN_1612; // @[CSR.scala 840:41]
  wire  _GEN_1613; // @[CSR.scala 838:89]
  wire [9:0] _T_671; // @[Cat.scala 29:58]
  wire [3:0] _T_675; // @[Cat.scala 29:58]
  wire [30:0] _T_676; // @[Cat.scala 29:58]
  wire [31:0] _T_678; // @[Cat.scala 29:58]
  wire [31:0] _T_680; // @[Cat.scala 29:58]
  wire [31:0] _T_682; // @[Cat.scala 29:58]
  wire [11:0] _T_692; // @[Cat.scala 29:58]
  wire [31:0] _T_693; // @[Cat.scala 29:58]
  wire [11:0] _T_703; // @[Cat.scala 29:58]
  wire [31:0] _T_704; // @[Cat.scala 29:58]
  wire [31:0] _T_707; // @[Cat.scala 29:58]
  wire [31:0] _T_710; // @[Cat.scala 29:58]
  wire [31:0] _T_713; // @[Cat.scala 29:58]
  wire [31:0] _T_716; // @[Cat.scala 29:58]
  wire [31:0] _T_727; // @[Cat.scala 29:58]
  wire [31:0] _T_729; // @[Cat.scala 29:58]
  wire [30:0] _T_734; // @[Cat.scala 29:58]
  wire [30:0] _T_739; // @[Cat.scala 29:58]
  wire [31:0] _T_742; // @[Cat.scala 29:58]
  wire [31:0] _T_745; // @[Cat.scala 29:58]
  wire [30:0] _T_748; // @[Cat.scala 29:58]
  wire [31:0] _T_751; // @[Cat.scala 29:58]
  wire [31:0] _GEN_1618; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1622; // @[Conditional.scala 39:67]
  wire  _GEN_1625; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1629; // @[Conditional.scala 39:67]
  wire  _GEN_1632; // @[Conditional.scala 39:67]
  wire  _GEN_1635; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1639; // @[Conditional.scala 39:67]
  wire  _GEN_1642; // @[Conditional.scala 39:67]
  wire  _GEN_1645; // @[Conditional.scala 39:67]
  wire  _GEN_1648; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1649; // @[Conditional.scala 39:67]
  wire  _GEN_1652; // @[Conditional.scala 39:67]
  wire  _GEN_1655; // @[Conditional.scala 39:67]
  wire  _GEN_1658; // @[Conditional.scala 39:67]
  wire  _GEN_1661; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1662; // @[Conditional.scala 39:67]
  wire  _GEN_1665; // @[Conditional.scala 39:67]
  wire  _GEN_1668; // @[Conditional.scala 39:67]
  wire  _GEN_1671; // @[Conditional.scala 39:67]
  wire  _GEN_1674; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1675; // @[Conditional.scala 39:67]
  wire  _GEN_1678; // @[Conditional.scala 39:67]
  wire  _GEN_1681; // @[Conditional.scala 39:67]
  wire  _GEN_1684; // @[Conditional.scala 39:67]
  wire  _GEN_1687; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1688; // @[Conditional.scala 39:67]
  wire  _GEN_1691; // @[Conditional.scala 39:67]
  wire  _GEN_1694; // @[Conditional.scala 39:67]
  wire  _GEN_1697; // @[Conditional.scala 39:67]
  wire  _GEN_1700; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1701; // @[Conditional.scala 39:67]
  wire  _GEN_1704; // @[Conditional.scala 39:67]
  wire  _GEN_1707; // @[Conditional.scala 39:67]
  wire  _GEN_1710; // @[Conditional.scala 39:67]
  wire  _GEN_1713; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1714; // @[Conditional.scala 39:67]
  wire  _GEN_1717; // @[Conditional.scala 39:67]
  wire  _GEN_1720; // @[Conditional.scala 39:67]
  wire  _GEN_1723; // @[Conditional.scala 39:67]
  wire  _GEN_1726; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1727; // @[Conditional.scala 39:67]
  wire  _GEN_1730; // @[Conditional.scala 39:67]
  wire  _GEN_1733; // @[Conditional.scala 39:67]
  wire  _GEN_1736; // @[Conditional.scala 39:67]
  wire  _GEN_1739; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1740; // @[Conditional.scala 39:67]
  wire  _GEN_1743; // @[Conditional.scala 39:67]
  wire  _GEN_1746; // @[Conditional.scala 39:67]
  wire  _GEN_1749; // @[Conditional.scala 39:67]
  wire  _GEN_1752; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1753; // @[Conditional.scala 39:67]
  wire  _GEN_1756; // @[Conditional.scala 39:67]
  wire  _GEN_1759; // @[Conditional.scala 39:67]
  wire  _GEN_1762; // @[Conditional.scala 39:67]
  wire  _GEN_1765; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1766; // @[Conditional.scala 39:67]
  wire  _GEN_1769; // @[Conditional.scala 39:67]
  wire  _GEN_1772; // @[Conditional.scala 39:67]
  wire  _GEN_1775; // @[Conditional.scala 39:67]
  wire  _GEN_1778; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1779; // @[Conditional.scala 39:67]
  wire  _GEN_1782; // @[Conditional.scala 39:67]
  wire  _GEN_1785; // @[Conditional.scala 39:67]
  wire  _GEN_1788; // @[Conditional.scala 39:67]
  wire  _GEN_1791; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1792; // @[Conditional.scala 39:67]
  wire  _GEN_1795; // @[Conditional.scala 39:67]
  wire  _GEN_1798; // @[Conditional.scala 39:67]
  wire  _GEN_1801; // @[Conditional.scala 39:67]
  wire  _GEN_1804; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1805; // @[Conditional.scala 39:67]
  wire  _GEN_1808; // @[Conditional.scala 39:67]
  wire  _GEN_1811; // @[Conditional.scala 39:67]
  wire  _GEN_1814; // @[Conditional.scala 39:67]
  wire  _GEN_1817; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1818; // @[Conditional.scala 39:67]
  wire  _GEN_1821; // @[Conditional.scala 39:67]
  wire  _GEN_1824; // @[Conditional.scala 39:67]
  wire  _GEN_1827; // @[Conditional.scala 39:67]
  wire  _GEN_1830; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1831; // @[Conditional.scala 39:67]
  wire  _GEN_1834; // @[Conditional.scala 39:67]
  wire  _GEN_1837; // @[Conditional.scala 39:67]
  wire  _GEN_1840; // @[Conditional.scala 39:67]
  wire  _GEN_1843; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1844; // @[Conditional.scala 39:67]
  wire  _GEN_1847; // @[Conditional.scala 39:67]
  wire  _GEN_1850; // @[Conditional.scala 39:67]
  wire  _GEN_1853; // @[Conditional.scala 39:67]
  wire  _GEN_1856; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1857; // @[Conditional.scala 39:67]
  wire  _GEN_1860; // @[Conditional.scala 39:67]
  wire  _GEN_1863; // @[Conditional.scala 39:67]
  wire  _GEN_1866; // @[Conditional.scala 39:67]
  wire  _GEN_1869; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1870; // @[Conditional.scala 39:67]
  wire  _GEN_1873; // @[Conditional.scala 39:67]
  wire  _GEN_1876; // @[Conditional.scala 39:67]
  wire  _GEN_1879; // @[Conditional.scala 39:67]
  wire  _GEN_1882; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1883; // @[Conditional.scala 39:67]
  wire  _GEN_1886; // @[Conditional.scala 39:67]
  wire  _GEN_1889; // @[Conditional.scala 39:67]
  wire  _GEN_1892; // @[Conditional.scala 39:67]
  wire  _GEN_1895; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1896; // @[Conditional.scala 39:67]
  wire  _GEN_1899; // @[Conditional.scala 39:67]
  wire  _GEN_1902; // @[Conditional.scala 39:67]
  wire  _GEN_1905; // @[Conditional.scala 39:67]
  wire  _GEN_1908; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1909; // @[Conditional.scala 39:67]
  wire  _GEN_1912; // @[Conditional.scala 39:67]
  wire  _GEN_1915; // @[Conditional.scala 39:67]
  wire  _GEN_1918; // @[Conditional.scala 39:67]
  wire  _GEN_1921; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1922; // @[Conditional.scala 39:67]
  wire  _GEN_1925; // @[Conditional.scala 39:67]
  wire  _GEN_1928; // @[Conditional.scala 39:67]
  wire  _GEN_1931; // @[Conditional.scala 39:67]
  wire  _GEN_1934; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1935; // @[Conditional.scala 39:67]
  wire  _GEN_1938; // @[Conditional.scala 39:67]
  wire  _GEN_1941; // @[Conditional.scala 39:67]
  wire  _GEN_1944; // @[Conditional.scala 39:67]
  wire  _GEN_1947; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1948; // @[Conditional.scala 39:67]
  wire  _GEN_1951; // @[Conditional.scala 39:67]
  wire  _GEN_1954; // @[Conditional.scala 39:67]
  wire  _GEN_1957; // @[Conditional.scala 39:67]
  wire  _GEN_1960; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1961; // @[Conditional.scala 39:67]
  wire  _GEN_1964; // @[Conditional.scala 39:67]
  wire  _GEN_1967; // @[Conditional.scala 39:67]
  wire  _GEN_1970; // @[Conditional.scala 39:67]
  wire  _GEN_1973; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1974; // @[Conditional.scala 39:67]
  wire  _GEN_1977; // @[Conditional.scala 39:67]
  wire  _GEN_1980; // @[Conditional.scala 39:67]
  wire  _GEN_1983; // @[Conditional.scala 39:67]
  wire  _GEN_1986; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_1987; // @[Conditional.scala 40:58]
  wire  _GEN_1990; // @[Conditional.scala 40:58]
  wire  _GEN_1993; // @[Conditional.scala 40:58]
  wire  _GEN_1996; // @[Conditional.scala 40:58]
  wire  _GEN_1999; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_2000; // @[CSR.scala 893:41]
  wire  _GEN_2003; // @[CSR.scala 893:41]
  wire  _GEN_2006; // @[CSR.scala 893:41]
  wire  _GEN_2009; // @[CSR.scala 893:41]
  wire  _GEN_2012; // @[CSR.scala 893:41]
  mmu_conv mmu_conv0 ( // @[CSR.scala 763:25]
    .io_rst_n(mmu_conv0_io_rst_n),
    .io_tlb0_vpn_i(mmu_conv0_io_tlb0_vpn_i),
    .io_tlb0_mask_i(mmu_conv0_io_tlb0_mask_i),
    .io_tlb0_pte_i(mmu_conv0_io_tlb0_pte_i),
    .io_tlb1_vpn_i(mmu_conv0_io_tlb1_vpn_i),
    .io_tlb1_mask_i(mmu_conv0_io_tlb1_mask_i),
    .io_tlb1_pte_i(mmu_conv0_io_tlb1_pte_i),
    .io_tlb2_vpn_i(mmu_conv0_io_tlb2_vpn_i),
    .io_tlb2_mask_i(mmu_conv0_io_tlb2_mask_i),
    .io_tlb2_pte_i(mmu_conv0_io_tlb2_pte_i),
    .io_tlb3_vpn_i(mmu_conv0_io_tlb3_vpn_i),
    .io_tlb3_mask_i(mmu_conv0_io_tlb3_mask_i),
    .io_tlb3_pte_i(mmu_conv0_io_tlb3_pte_i),
    .io_tlb4_vpn_i(mmu_conv0_io_tlb4_vpn_i),
    .io_tlb4_mask_i(mmu_conv0_io_tlb4_mask_i),
    .io_tlb4_pte_i(mmu_conv0_io_tlb4_pte_i),
    .io_tlb5_vpn_i(mmu_conv0_io_tlb5_vpn_i),
    .io_tlb5_mask_i(mmu_conv0_io_tlb5_mask_i),
    .io_tlb5_pte_i(mmu_conv0_io_tlb5_pte_i),
    .io_tlb6_vpn_i(mmu_conv0_io_tlb6_vpn_i),
    .io_tlb6_mask_i(mmu_conv0_io_tlb6_mask_i),
    .io_tlb6_pte_i(mmu_conv0_io_tlb6_pte_i),
    .io_tlb7_vpn_i(mmu_conv0_io_tlb7_vpn_i),
    .io_tlb7_mask_i(mmu_conv0_io_tlb7_mask_i),
    .io_tlb7_pte_i(mmu_conv0_io_tlb7_pte_i),
    .io_tlb8_vpn_i(mmu_conv0_io_tlb8_vpn_i),
    .io_tlb8_mask_i(mmu_conv0_io_tlb8_mask_i),
    .io_tlb8_pte_i(mmu_conv0_io_tlb8_pte_i),
    .io_tlb9_vpn_i(mmu_conv0_io_tlb9_vpn_i),
    .io_tlb9_mask_i(mmu_conv0_io_tlb9_mask_i),
    .io_tlb9_pte_i(mmu_conv0_io_tlb9_pte_i),
    .io_tlb10_vpn_i(mmu_conv0_io_tlb10_vpn_i),
    .io_tlb10_mask_i(mmu_conv0_io_tlb10_mask_i),
    .io_tlb10_pte_i(mmu_conv0_io_tlb10_pte_i),
    .io_tlb11_vpn_i(mmu_conv0_io_tlb11_vpn_i),
    .io_tlb11_mask_i(mmu_conv0_io_tlb11_mask_i),
    .io_tlb11_pte_i(mmu_conv0_io_tlb11_pte_i),
    .io_tlb12_vpn_i(mmu_conv0_io_tlb12_vpn_i),
    .io_tlb12_mask_i(mmu_conv0_io_tlb12_mask_i),
    .io_tlb12_pte_i(mmu_conv0_io_tlb12_pte_i),
    .io_tlb13_vpn_i(mmu_conv0_io_tlb13_vpn_i),
    .io_tlb13_mask_i(mmu_conv0_io_tlb13_mask_i),
    .io_tlb13_pte_i(mmu_conv0_io_tlb13_pte_i),
    .io_tlb14_vpn_i(mmu_conv0_io_tlb14_vpn_i),
    .io_tlb14_mask_i(mmu_conv0_io_tlb14_mask_i),
    .io_tlb14_pte_i(mmu_conv0_io_tlb14_pte_i),
    .io_tlb15_vpn_i(mmu_conv0_io_tlb15_vpn_i),
    .io_tlb15_mask_i(mmu_conv0_io_tlb15_mask_i),
    .io_tlb15_pte_i(mmu_conv0_io_tlb15_pte_i),
    .io_vm_i(mmu_conv0_io_vm_i),
    .io_prv_i(mmu_conv0_io_prv_i),
    .io_mxr_i(mmu_conv0_io_mxr_i),
    .io_ce_i(mmu_conv0_io_ce_i),
    .io_ex_i(mmu_conv0_io_ex_i),
    .io_we_i(mmu_conv0_io_we_i),
    .io_vir_addr_i(mmu_conv0_io_vir_addr_i),
    .io_phy_addr_o(mmu_conv0_io_phy_addr_o),
    .io_tlb_exception_o(mmu_conv0_io_tlb_exception_o),
    .io_tlb_update_o(mmu_conv0_io_tlb_update_o),
    .io_hit_index_o(mmu_conv0_io_hit_index_o)
  );
  mmu_conv mmu_conv1 ( // @[CSR.scala 799:25]
    .io_rst_n(mmu_conv1_io_rst_n),
    .io_tlb0_vpn_i(mmu_conv1_io_tlb0_vpn_i),
    .io_tlb0_mask_i(mmu_conv1_io_tlb0_mask_i),
    .io_tlb0_pte_i(mmu_conv1_io_tlb0_pte_i),
    .io_tlb1_vpn_i(mmu_conv1_io_tlb1_vpn_i),
    .io_tlb1_mask_i(mmu_conv1_io_tlb1_mask_i),
    .io_tlb1_pte_i(mmu_conv1_io_tlb1_pte_i),
    .io_tlb2_vpn_i(mmu_conv1_io_tlb2_vpn_i),
    .io_tlb2_mask_i(mmu_conv1_io_tlb2_mask_i),
    .io_tlb2_pte_i(mmu_conv1_io_tlb2_pte_i),
    .io_tlb3_vpn_i(mmu_conv1_io_tlb3_vpn_i),
    .io_tlb3_mask_i(mmu_conv1_io_tlb3_mask_i),
    .io_tlb3_pte_i(mmu_conv1_io_tlb3_pte_i),
    .io_tlb4_vpn_i(mmu_conv1_io_tlb4_vpn_i),
    .io_tlb4_mask_i(mmu_conv1_io_tlb4_mask_i),
    .io_tlb4_pte_i(mmu_conv1_io_tlb4_pte_i),
    .io_tlb5_vpn_i(mmu_conv1_io_tlb5_vpn_i),
    .io_tlb5_mask_i(mmu_conv1_io_tlb5_mask_i),
    .io_tlb5_pte_i(mmu_conv1_io_tlb5_pte_i),
    .io_tlb6_vpn_i(mmu_conv1_io_tlb6_vpn_i),
    .io_tlb6_mask_i(mmu_conv1_io_tlb6_mask_i),
    .io_tlb6_pte_i(mmu_conv1_io_tlb6_pte_i),
    .io_tlb7_vpn_i(mmu_conv1_io_tlb7_vpn_i),
    .io_tlb7_mask_i(mmu_conv1_io_tlb7_mask_i),
    .io_tlb7_pte_i(mmu_conv1_io_tlb7_pte_i),
    .io_tlb8_vpn_i(mmu_conv1_io_tlb8_vpn_i),
    .io_tlb8_mask_i(mmu_conv1_io_tlb8_mask_i),
    .io_tlb8_pte_i(mmu_conv1_io_tlb8_pte_i),
    .io_tlb9_vpn_i(mmu_conv1_io_tlb9_vpn_i),
    .io_tlb9_mask_i(mmu_conv1_io_tlb9_mask_i),
    .io_tlb9_pte_i(mmu_conv1_io_tlb9_pte_i),
    .io_tlb10_vpn_i(mmu_conv1_io_tlb10_vpn_i),
    .io_tlb10_mask_i(mmu_conv1_io_tlb10_mask_i),
    .io_tlb10_pte_i(mmu_conv1_io_tlb10_pte_i),
    .io_tlb11_vpn_i(mmu_conv1_io_tlb11_vpn_i),
    .io_tlb11_mask_i(mmu_conv1_io_tlb11_mask_i),
    .io_tlb11_pte_i(mmu_conv1_io_tlb11_pte_i),
    .io_tlb12_vpn_i(mmu_conv1_io_tlb12_vpn_i),
    .io_tlb12_mask_i(mmu_conv1_io_tlb12_mask_i),
    .io_tlb12_pte_i(mmu_conv1_io_tlb12_pte_i),
    .io_tlb13_vpn_i(mmu_conv1_io_tlb13_vpn_i),
    .io_tlb13_mask_i(mmu_conv1_io_tlb13_mask_i),
    .io_tlb13_pte_i(mmu_conv1_io_tlb13_pte_i),
    .io_tlb14_vpn_i(mmu_conv1_io_tlb14_vpn_i),
    .io_tlb14_mask_i(mmu_conv1_io_tlb14_mask_i),
    .io_tlb14_pte_i(mmu_conv1_io_tlb14_pte_i),
    .io_tlb15_vpn_i(mmu_conv1_io_tlb15_vpn_i),
    .io_tlb15_mask_i(mmu_conv1_io_tlb15_mask_i),
    .io_tlb15_pte_i(mmu_conv1_io_tlb15_pte_i),
    .io_vm_i(mmu_conv1_io_vm_i),
    .io_prv_i(mmu_conv1_io_prv_i),
    .io_mxr_i(mmu_conv1_io_mxr_i),
    .io_ce_i(mmu_conv1_io_ce_i),
    .io_ex_i(mmu_conv1_io_ex_i),
    .io_we_i(mmu_conv1_io_we_i),
    .io_vir_addr_i(mmu_conv1_io_vir_addr_i),
    .io_phy_addr_o(mmu_conv1_io_phy_addr_o),
    .io_tlb_exception_o(mmu_conv1_io_tlb_exception_o),
    .io_tlb_update_o(mmu_conv1_io_tlb_update_o),
    .io_hit_index_o(mmu_conv1_io_hit_index_o)
  );
  assign mtlbvpn__T_480_addr = 4'h0;
  assign mtlbvpn__T_480_data = mtlbvpn[mtlbvpn__T_480_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_483_addr = 4'h1;
  assign mtlbvpn__T_483_data = mtlbvpn[mtlbvpn__T_483_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_486_addr = 4'h2;
  assign mtlbvpn__T_486_data = mtlbvpn[mtlbvpn__T_486_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_489_addr = 4'h3;
  assign mtlbvpn__T_489_data = mtlbvpn[mtlbvpn__T_489_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_492_addr = 4'h4;
  assign mtlbvpn__T_492_data = mtlbvpn[mtlbvpn__T_492_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_495_addr = 4'h5;
  assign mtlbvpn__T_495_data = mtlbvpn[mtlbvpn__T_495_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_498_addr = 4'h6;
  assign mtlbvpn__T_498_data = mtlbvpn[mtlbvpn__T_498_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_501_addr = 4'h7;
  assign mtlbvpn__T_501_data = mtlbvpn[mtlbvpn__T_501_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_504_addr = 4'h8;
  assign mtlbvpn__T_504_data = mtlbvpn[mtlbvpn__T_504_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_507_addr = 4'h9;
  assign mtlbvpn__T_507_data = mtlbvpn[mtlbvpn__T_507_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_510_addr = 4'ha;
  assign mtlbvpn__T_510_data = mtlbvpn[mtlbvpn__T_510_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_513_addr = 4'hb;
  assign mtlbvpn__T_513_data = mtlbvpn[mtlbvpn__T_513_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_516_addr = 4'hc;
  assign mtlbvpn__T_516_data = mtlbvpn[mtlbvpn__T_516_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_519_addr = 4'hd;
  assign mtlbvpn__T_519_data = mtlbvpn[mtlbvpn__T_519_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_522_addr = 4'he;
  assign mtlbvpn__T_522_data = mtlbvpn[mtlbvpn__T_522_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_525_addr = 4'hf;
  assign mtlbvpn__T_525_data = mtlbvpn[mtlbvpn__T_525_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_528_addr = 4'h0;
  assign mtlbvpn__T_528_data = mtlbvpn[mtlbvpn__T_528_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_531_addr = 4'h1;
  assign mtlbvpn__T_531_data = mtlbvpn[mtlbvpn__T_531_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_534_addr = 4'h2;
  assign mtlbvpn__T_534_data = mtlbvpn[mtlbvpn__T_534_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_537_addr = 4'h3;
  assign mtlbvpn__T_537_data = mtlbvpn[mtlbvpn__T_537_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_540_addr = 4'h4;
  assign mtlbvpn__T_540_data = mtlbvpn[mtlbvpn__T_540_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_543_addr = 4'h5;
  assign mtlbvpn__T_543_data = mtlbvpn[mtlbvpn__T_543_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_546_addr = 4'h6;
  assign mtlbvpn__T_546_data = mtlbvpn[mtlbvpn__T_546_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_549_addr = 4'h7;
  assign mtlbvpn__T_549_data = mtlbvpn[mtlbvpn__T_549_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_552_addr = 4'h8;
  assign mtlbvpn__T_552_data = mtlbvpn[mtlbvpn__T_552_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_555_addr = 4'h9;
  assign mtlbvpn__T_555_data = mtlbvpn[mtlbvpn__T_555_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_558_addr = 4'ha;
  assign mtlbvpn__T_558_data = mtlbvpn[mtlbvpn__T_558_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_561_addr = 4'hb;
  assign mtlbvpn__T_561_data = mtlbvpn[mtlbvpn__T_561_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_564_addr = 4'hc;
  assign mtlbvpn__T_564_data = mtlbvpn[mtlbvpn__T_564_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_567_addr = 4'hd;
  assign mtlbvpn__T_567_data = mtlbvpn[mtlbvpn__T_567_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_570_addr = 4'he;
  assign mtlbvpn__T_570_data = mtlbvpn[mtlbvpn__T_570_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_573_addr = 4'hf;
  assign mtlbvpn__T_573_data = mtlbvpn[mtlbvpn__T_573_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_753_addr = mtlbindex;
  assign mtlbvpn__T_753_data = mtlbvpn[mtlbvpn__T_753_addr]; // @[CSR.scala 121:26]
  assign mtlbvpn__T_192_data = 32'h0;
  assign mtlbvpn__T_192_addr = 4'h0;
  assign mtlbvpn__T_192_mask = 1'h1;
  assign mtlbvpn__T_192_en = ~io_rst_n;
  assign mtlbvpn__T_196_data = 32'h0;
  assign mtlbvpn__T_196_addr = 4'h1;
  assign mtlbvpn__T_196_mask = 1'h1;
  assign mtlbvpn__T_196_en = ~io_rst_n;
  assign mtlbvpn__T_200_data = 32'h0;
  assign mtlbvpn__T_200_addr = 4'h2;
  assign mtlbvpn__T_200_mask = 1'h1;
  assign mtlbvpn__T_200_en = ~io_rst_n;
  assign mtlbvpn__T_204_data = 32'h0;
  assign mtlbvpn__T_204_addr = 4'h3;
  assign mtlbvpn__T_204_mask = 1'h1;
  assign mtlbvpn__T_204_en = ~io_rst_n;
  assign mtlbvpn__T_208_data = 32'h0;
  assign mtlbvpn__T_208_addr = 4'h4;
  assign mtlbvpn__T_208_mask = 1'h1;
  assign mtlbvpn__T_208_en = ~io_rst_n;
  assign mtlbvpn__T_212_data = 32'h0;
  assign mtlbvpn__T_212_addr = 4'h5;
  assign mtlbvpn__T_212_mask = 1'h1;
  assign mtlbvpn__T_212_en = ~io_rst_n;
  assign mtlbvpn__T_216_data = 32'h0;
  assign mtlbvpn__T_216_addr = 4'h6;
  assign mtlbvpn__T_216_mask = 1'h1;
  assign mtlbvpn__T_216_en = ~io_rst_n;
  assign mtlbvpn__T_220_data = 32'h0;
  assign mtlbvpn__T_220_addr = 4'h7;
  assign mtlbvpn__T_220_mask = 1'h1;
  assign mtlbvpn__T_220_en = ~io_rst_n;
  assign mtlbvpn__T_224_data = 32'h0;
  assign mtlbvpn__T_224_addr = 4'h8;
  assign mtlbvpn__T_224_mask = 1'h1;
  assign mtlbvpn__T_224_en = ~io_rst_n;
  assign mtlbvpn__T_228_data = 32'h0;
  assign mtlbvpn__T_228_addr = 4'h9;
  assign mtlbvpn__T_228_mask = 1'h1;
  assign mtlbvpn__T_228_en = ~io_rst_n;
  assign mtlbvpn__T_232_data = 32'h0;
  assign mtlbvpn__T_232_addr = 4'ha;
  assign mtlbvpn__T_232_mask = 1'h1;
  assign mtlbvpn__T_232_en = ~io_rst_n;
  assign mtlbvpn__T_236_data = 32'h0;
  assign mtlbvpn__T_236_addr = 4'hb;
  assign mtlbvpn__T_236_mask = 1'h1;
  assign mtlbvpn__T_236_en = ~io_rst_n;
  assign mtlbvpn__T_240_data = 32'h0;
  assign mtlbvpn__T_240_addr = 4'hc;
  assign mtlbvpn__T_240_mask = 1'h1;
  assign mtlbvpn__T_240_en = ~io_rst_n;
  assign mtlbvpn__T_244_data = 32'h0;
  assign mtlbvpn__T_244_addr = 4'hd;
  assign mtlbvpn__T_244_mask = 1'h1;
  assign mtlbvpn__T_244_en = ~io_rst_n;
  assign mtlbvpn__T_248_data = 32'h0;
  assign mtlbvpn__T_248_addr = 4'he;
  assign mtlbvpn__T_248_mask = 1'h1;
  assign mtlbvpn__T_248_en = ~io_rst_n;
  assign mtlbvpn__T_252_data = 32'h0;
  assign mtlbvpn__T_252_addr = 4'hf;
  assign mtlbvpn__T_252_mask = 1'h1;
  assign mtlbvpn__T_252_en = ~io_rst_n;
  assign mtlbvpn__T_469_data = io_data_i;
  assign mtlbvpn__T_469_addr = mtlbindex;
  assign mtlbvpn__T_469_mask = 1'h1;
  assign mtlbvpn__T_469_en = io_rst_n ? _GEN_1509 : 1'h0;
  assign mtlbmask__T_482_addr = 4'h0;
  assign mtlbmask__T_482_data = mtlbmask[mtlbmask__T_482_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_485_addr = 4'h1;
  assign mtlbmask__T_485_data = mtlbmask[mtlbmask__T_485_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_488_addr = 4'h2;
  assign mtlbmask__T_488_data = mtlbmask[mtlbmask__T_488_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_491_addr = 4'h3;
  assign mtlbmask__T_491_data = mtlbmask[mtlbmask__T_491_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_494_addr = 4'h4;
  assign mtlbmask__T_494_data = mtlbmask[mtlbmask__T_494_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_497_addr = 4'h5;
  assign mtlbmask__T_497_data = mtlbmask[mtlbmask__T_497_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_500_addr = 4'h6;
  assign mtlbmask__T_500_data = mtlbmask[mtlbmask__T_500_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_503_addr = 4'h7;
  assign mtlbmask__T_503_data = mtlbmask[mtlbmask__T_503_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_506_addr = 4'h8;
  assign mtlbmask__T_506_data = mtlbmask[mtlbmask__T_506_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_509_addr = 4'h9;
  assign mtlbmask__T_509_data = mtlbmask[mtlbmask__T_509_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_512_addr = 4'ha;
  assign mtlbmask__T_512_data = mtlbmask[mtlbmask__T_512_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_515_addr = 4'hb;
  assign mtlbmask__T_515_data = mtlbmask[mtlbmask__T_515_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_518_addr = 4'hc;
  assign mtlbmask__T_518_data = mtlbmask[mtlbmask__T_518_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_521_addr = 4'hd;
  assign mtlbmask__T_521_data = mtlbmask[mtlbmask__T_521_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_524_addr = 4'he;
  assign mtlbmask__T_524_data = mtlbmask[mtlbmask__T_524_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_527_addr = 4'hf;
  assign mtlbmask__T_527_data = mtlbmask[mtlbmask__T_527_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_530_addr = 4'h0;
  assign mtlbmask__T_530_data = mtlbmask[mtlbmask__T_530_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_533_addr = 4'h1;
  assign mtlbmask__T_533_data = mtlbmask[mtlbmask__T_533_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_536_addr = 4'h2;
  assign mtlbmask__T_536_data = mtlbmask[mtlbmask__T_536_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_539_addr = 4'h3;
  assign mtlbmask__T_539_data = mtlbmask[mtlbmask__T_539_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_542_addr = 4'h4;
  assign mtlbmask__T_542_data = mtlbmask[mtlbmask__T_542_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_545_addr = 4'h5;
  assign mtlbmask__T_545_data = mtlbmask[mtlbmask__T_545_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_548_addr = 4'h6;
  assign mtlbmask__T_548_data = mtlbmask[mtlbmask__T_548_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_551_addr = 4'h7;
  assign mtlbmask__T_551_data = mtlbmask[mtlbmask__T_551_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_554_addr = 4'h8;
  assign mtlbmask__T_554_data = mtlbmask[mtlbmask__T_554_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_557_addr = 4'h9;
  assign mtlbmask__T_557_data = mtlbmask[mtlbmask__T_557_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_560_addr = 4'ha;
  assign mtlbmask__T_560_data = mtlbmask[mtlbmask__T_560_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_563_addr = 4'hb;
  assign mtlbmask__T_563_data = mtlbmask[mtlbmask__T_563_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_566_addr = 4'hc;
  assign mtlbmask__T_566_data = mtlbmask[mtlbmask__T_566_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_569_addr = 4'hd;
  assign mtlbmask__T_569_data = mtlbmask[mtlbmask__T_569_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_572_addr = 4'he;
  assign mtlbmask__T_572_data = mtlbmask[mtlbmask__T_572_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_575_addr = 4'hf;
  assign mtlbmask__T_575_data = mtlbmask[mtlbmask__T_575_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_755_addr = mtlbindex;
  assign mtlbmask__T_755_data = mtlbmask[mtlbmask__T_755_addr]; // @[CSR.scala 122:26]
  assign mtlbmask__T_193_data = 32'h0;
  assign mtlbmask__T_193_addr = 4'h0;
  assign mtlbmask__T_193_mask = 1'h1;
  assign mtlbmask__T_193_en = ~io_rst_n;
  assign mtlbmask__T_197_data = 32'h0;
  assign mtlbmask__T_197_addr = 4'h1;
  assign mtlbmask__T_197_mask = 1'h1;
  assign mtlbmask__T_197_en = ~io_rst_n;
  assign mtlbmask__T_201_data = 32'h0;
  assign mtlbmask__T_201_addr = 4'h2;
  assign mtlbmask__T_201_mask = 1'h1;
  assign mtlbmask__T_201_en = ~io_rst_n;
  assign mtlbmask__T_205_data = 32'h0;
  assign mtlbmask__T_205_addr = 4'h3;
  assign mtlbmask__T_205_mask = 1'h1;
  assign mtlbmask__T_205_en = ~io_rst_n;
  assign mtlbmask__T_209_data = 32'h0;
  assign mtlbmask__T_209_addr = 4'h4;
  assign mtlbmask__T_209_mask = 1'h1;
  assign mtlbmask__T_209_en = ~io_rst_n;
  assign mtlbmask__T_213_data = 32'h0;
  assign mtlbmask__T_213_addr = 4'h5;
  assign mtlbmask__T_213_mask = 1'h1;
  assign mtlbmask__T_213_en = ~io_rst_n;
  assign mtlbmask__T_217_data = 32'h0;
  assign mtlbmask__T_217_addr = 4'h6;
  assign mtlbmask__T_217_mask = 1'h1;
  assign mtlbmask__T_217_en = ~io_rst_n;
  assign mtlbmask__T_221_data = 32'h0;
  assign mtlbmask__T_221_addr = 4'h7;
  assign mtlbmask__T_221_mask = 1'h1;
  assign mtlbmask__T_221_en = ~io_rst_n;
  assign mtlbmask__T_225_data = 32'h0;
  assign mtlbmask__T_225_addr = 4'h8;
  assign mtlbmask__T_225_mask = 1'h1;
  assign mtlbmask__T_225_en = ~io_rst_n;
  assign mtlbmask__T_229_data = 32'h0;
  assign mtlbmask__T_229_addr = 4'h9;
  assign mtlbmask__T_229_mask = 1'h1;
  assign mtlbmask__T_229_en = ~io_rst_n;
  assign mtlbmask__T_233_data = 32'h0;
  assign mtlbmask__T_233_addr = 4'ha;
  assign mtlbmask__T_233_mask = 1'h1;
  assign mtlbmask__T_233_en = ~io_rst_n;
  assign mtlbmask__T_237_data = 32'h0;
  assign mtlbmask__T_237_addr = 4'hb;
  assign mtlbmask__T_237_mask = 1'h1;
  assign mtlbmask__T_237_en = ~io_rst_n;
  assign mtlbmask__T_241_data = 32'h0;
  assign mtlbmask__T_241_addr = 4'hc;
  assign mtlbmask__T_241_mask = 1'h1;
  assign mtlbmask__T_241_en = ~io_rst_n;
  assign mtlbmask__T_245_data = 32'h0;
  assign mtlbmask__T_245_addr = 4'hd;
  assign mtlbmask__T_245_mask = 1'h1;
  assign mtlbmask__T_245_en = ~io_rst_n;
  assign mtlbmask__T_249_data = 32'h0;
  assign mtlbmask__T_249_addr = 4'he;
  assign mtlbmask__T_249_mask = 1'h1;
  assign mtlbmask__T_249_en = ~io_rst_n;
  assign mtlbmask__T_253_data = 32'h0;
  assign mtlbmask__T_253_addr = 4'hf;
  assign mtlbmask__T_253_mask = 1'h1;
  assign mtlbmask__T_253_en = ~io_rst_n;
  assign mtlbmask__T_471_data = io_data_i;
  assign mtlbmask__T_471_addr = mtlbindex;
  assign mtlbmask__T_471_mask = 1'h1;
  assign mtlbmask__T_471_en = io_rst_n ? _GEN_1514 : 1'h0;
  assign mtlbpte__T_481_addr = 4'h0;
  assign mtlbpte__T_481_data = mtlbpte[mtlbpte__T_481_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_484_addr = 4'h1;
  assign mtlbpte__T_484_data = mtlbpte[mtlbpte__T_484_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_487_addr = 4'h2;
  assign mtlbpte__T_487_data = mtlbpte[mtlbpte__T_487_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_490_addr = 4'h3;
  assign mtlbpte__T_490_data = mtlbpte[mtlbpte__T_490_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_493_addr = 4'h4;
  assign mtlbpte__T_493_data = mtlbpte[mtlbpte__T_493_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_496_addr = 4'h5;
  assign mtlbpte__T_496_data = mtlbpte[mtlbpte__T_496_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_499_addr = 4'h6;
  assign mtlbpte__T_499_data = mtlbpte[mtlbpte__T_499_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_502_addr = 4'h7;
  assign mtlbpte__T_502_data = mtlbpte[mtlbpte__T_502_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_505_addr = 4'h8;
  assign mtlbpte__T_505_data = mtlbpte[mtlbpte__T_505_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_508_addr = 4'h9;
  assign mtlbpte__T_508_data = mtlbpte[mtlbpte__T_508_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_511_addr = 4'ha;
  assign mtlbpte__T_511_data = mtlbpte[mtlbpte__T_511_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_514_addr = 4'hb;
  assign mtlbpte__T_514_data = mtlbpte[mtlbpte__T_514_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_517_addr = 4'hc;
  assign mtlbpte__T_517_data = mtlbpte[mtlbpte__T_517_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_520_addr = 4'hd;
  assign mtlbpte__T_520_data = mtlbpte[mtlbpte__T_520_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_523_addr = 4'he;
  assign mtlbpte__T_523_data = mtlbpte[mtlbpte__T_523_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_526_addr = 4'hf;
  assign mtlbpte__T_526_data = mtlbpte[mtlbpte__T_526_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_529_addr = 4'h0;
  assign mtlbpte__T_529_data = mtlbpte[mtlbpte__T_529_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_532_addr = 4'h1;
  assign mtlbpte__T_532_data = mtlbpte[mtlbpte__T_532_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_535_addr = 4'h2;
  assign mtlbpte__T_535_data = mtlbpte[mtlbpte__T_535_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_538_addr = 4'h3;
  assign mtlbpte__T_538_data = mtlbpte[mtlbpte__T_538_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_541_addr = 4'h4;
  assign mtlbpte__T_541_data = mtlbpte[mtlbpte__T_541_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_544_addr = 4'h5;
  assign mtlbpte__T_544_data = mtlbpte[mtlbpte__T_544_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_547_addr = 4'h6;
  assign mtlbpte__T_547_data = mtlbpte[mtlbpte__T_547_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_550_addr = 4'h7;
  assign mtlbpte__T_550_data = mtlbpte[mtlbpte__T_550_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_553_addr = 4'h8;
  assign mtlbpte__T_553_data = mtlbpte[mtlbpte__T_553_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_556_addr = 4'h9;
  assign mtlbpte__T_556_data = mtlbpte[mtlbpte__T_556_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_559_addr = 4'ha;
  assign mtlbpte__T_559_data = mtlbpte[mtlbpte__T_559_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_562_addr = 4'hb;
  assign mtlbpte__T_562_data = mtlbpte[mtlbpte__T_562_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_565_addr = 4'hc;
  assign mtlbpte__T_565_data = mtlbpte[mtlbpte__T_565_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_568_addr = 4'hd;
  assign mtlbpte__T_568_data = mtlbpte[mtlbpte__T_568_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_571_addr = 4'he;
  assign mtlbpte__T_571_data = mtlbpte[mtlbpte__T_571_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_574_addr = 4'hf;
  assign mtlbpte__T_574_data = mtlbpte[mtlbpte__T_574_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_757_addr = mtlbindex;
  assign mtlbpte__T_757_data = mtlbpte[mtlbpte__T_757_addr]; // @[CSR.scala 123:26]
  assign mtlbpte__T_194_data = 32'h0;
  assign mtlbpte__T_194_addr = 4'h0;
  assign mtlbpte__T_194_mask = 1'h1;
  assign mtlbpte__T_194_en = ~io_rst_n;
  assign mtlbpte__T_198_data = 32'h0;
  assign mtlbpte__T_198_addr = 4'h1;
  assign mtlbpte__T_198_mask = 1'h1;
  assign mtlbpte__T_198_en = ~io_rst_n;
  assign mtlbpte__T_202_data = 32'h0;
  assign mtlbpte__T_202_addr = 4'h2;
  assign mtlbpte__T_202_mask = 1'h1;
  assign mtlbpte__T_202_en = ~io_rst_n;
  assign mtlbpte__T_206_data = 32'h0;
  assign mtlbpte__T_206_addr = 4'h3;
  assign mtlbpte__T_206_mask = 1'h1;
  assign mtlbpte__T_206_en = ~io_rst_n;
  assign mtlbpte__T_210_data = 32'h0;
  assign mtlbpte__T_210_addr = 4'h4;
  assign mtlbpte__T_210_mask = 1'h1;
  assign mtlbpte__T_210_en = ~io_rst_n;
  assign mtlbpte__T_214_data = 32'h0;
  assign mtlbpte__T_214_addr = 4'h5;
  assign mtlbpte__T_214_mask = 1'h1;
  assign mtlbpte__T_214_en = ~io_rst_n;
  assign mtlbpte__T_218_data = 32'h0;
  assign mtlbpte__T_218_addr = 4'h6;
  assign mtlbpte__T_218_mask = 1'h1;
  assign mtlbpte__T_218_en = ~io_rst_n;
  assign mtlbpte__T_222_data = 32'h0;
  assign mtlbpte__T_222_addr = 4'h7;
  assign mtlbpte__T_222_mask = 1'h1;
  assign mtlbpte__T_222_en = ~io_rst_n;
  assign mtlbpte__T_226_data = 32'h0;
  assign mtlbpte__T_226_addr = 4'h8;
  assign mtlbpte__T_226_mask = 1'h1;
  assign mtlbpte__T_226_en = ~io_rst_n;
  assign mtlbpte__T_230_data = 32'h0;
  assign mtlbpte__T_230_addr = 4'h9;
  assign mtlbpte__T_230_mask = 1'h1;
  assign mtlbpte__T_230_en = ~io_rst_n;
  assign mtlbpte__T_234_data = 32'h0;
  assign mtlbpte__T_234_addr = 4'ha;
  assign mtlbpte__T_234_mask = 1'h1;
  assign mtlbpte__T_234_en = ~io_rst_n;
  assign mtlbpte__T_238_data = 32'h0;
  assign mtlbpte__T_238_addr = 4'hb;
  assign mtlbpte__T_238_mask = 1'h1;
  assign mtlbpte__T_238_en = ~io_rst_n;
  assign mtlbpte__T_242_data = 32'h0;
  assign mtlbpte__T_242_addr = 4'hc;
  assign mtlbpte__T_242_mask = 1'h1;
  assign mtlbpte__T_242_en = ~io_rst_n;
  assign mtlbpte__T_246_data = 32'h0;
  assign mtlbpte__T_246_addr = 4'hd;
  assign mtlbpte__T_246_mask = 1'h1;
  assign mtlbpte__T_246_en = ~io_rst_n;
  assign mtlbpte__T_250_data = 32'h0;
  assign mtlbpte__T_250_addr = 4'he;
  assign mtlbpte__T_250_mask = 1'h1;
  assign mtlbpte__T_250_en = ~io_rst_n;
  assign mtlbpte__T_254_data = 32'h0;
  assign mtlbpte__T_254_addr = 4'hf;
  assign mtlbpte__T_254_mask = 1'h1;
  assign mtlbpte__T_254_en = ~io_rst_n;
  assign mtlbpte__T_473_data = io_data_i;
  assign mtlbpte__T_473_addr = mtlbindex;
  assign mtlbpte__T_473_mask = 1'h1;
  assign mtlbpte__T_473_en = io_rst_n ? _GEN_1519 : 1'h0;
  assign mtlbptevaddr__T_759_addr = mtlbindex;
  assign mtlbptevaddr__T_759_data = mtlbptevaddr[mtlbptevaddr__T_759_addr]; // @[CSR.scala 124:26]
  assign mtlbptevaddr__T_195_data = 32'h0;
  assign mtlbptevaddr__T_195_addr = 4'h0;
  assign mtlbptevaddr__T_195_mask = 1'h1;
  assign mtlbptevaddr__T_195_en = ~io_rst_n;
  assign mtlbptevaddr__T_199_data = 32'h0;
  assign mtlbptevaddr__T_199_addr = 4'h1;
  assign mtlbptevaddr__T_199_mask = 1'h1;
  assign mtlbptevaddr__T_199_en = ~io_rst_n;
  assign mtlbptevaddr__T_203_data = 32'h0;
  assign mtlbptevaddr__T_203_addr = 4'h2;
  assign mtlbptevaddr__T_203_mask = 1'h1;
  assign mtlbptevaddr__T_203_en = ~io_rst_n;
  assign mtlbptevaddr__T_207_data = 32'h0;
  assign mtlbptevaddr__T_207_addr = 4'h3;
  assign mtlbptevaddr__T_207_mask = 1'h1;
  assign mtlbptevaddr__T_207_en = ~io_rst_n;
  assign mtlbptevaddr__T_211_data = 32'h0;
  assign mtlbptevaddr__T_211_addr = 4'h4;
  assign mtlbptevaddr__T_211_mask = 1'h1;
  assign mtlbptevaddr__T_211_en = ~io_rst_n;
  assign mtlbptevaddr__T_215_data = 32'h0;
  assign mtlbptevaddr__T_215_addr = 4'h5;
  assign mtlbptevaddr__T_215_mask = 1'h1;
  assign mtlbptevaddr__T_215_en = ~io_rst_n;
  assign mtlbptevaddr__T_219_data = 32'h0;
  assign mtlbptevaddr__T_219_addr = 4'h6;
  assign mtlbptevaddr__T_219_mask = 1'h1;
  assign mtlbptevaddr__T_219_en = ~io_rst_n;
  assign mtlbptevaddr__T_223_data = 32'h0;
  assign mtlbptevaddr__T_223_addr = 4'h7;
  assign mtlbptevaddr__T_223_mask = 1'h1;
  assign mtlbptevaddr__T_223_en = ~io_rst_n;
  assign mtlbptevaddr__T_227_data = 32'h0;
  assign mtlbptevaddr__T_227_addr = 4'h8;
  assign mtlbptevaddr__T_227_mask = 1'h1;
  assign mtlbptevaddr__T_227_en = ~io_rst_n;
  assign mtlbptevaddr__T_231_data = 32'h0;
  assign mtlbptevaddr__T_231_addr = 4'h9;
  assign mtlbptevaddr__T_231_mask = 1'h1;
  assign mtlbptevaddr__T_231_en = ~io_rst_n;
  assign mtlbptevaddr__T_235_data = 32'h0;
  assign mtlbptevaddr__T_235_addr = 4'ha;
  assign mtlbptevaddr__T_235_mask = 1'h1;
  assign mtlbptevaddr__T_235_en = ~io_rst_n;
  assign mtlbptevaddr__T_239_data = 32'h0;
  assign mtlbptevaddr__T_239_addr = 4'hb;
  assign mtlbptevaddr__T_239_mask = 1'h1;
  assign mtlbptevaddr__T_239_en = ~io_rst_n;
  assign mtlbptevaddr__T_243_data = 32'h0;
  assign mtlbptevaddr__T_243_addr = 4'hc;
  assign mtlbptevaddr__T_243_mask = 1'h1;
  assign mtlbptevaddr__T_243_en = ~io_rst_n;
  assign mtlbptevaddr__T_247_data = 32'h0;
  assign mtlbptevaddr__T_247_addr = 4'hd;
  assign mtlbptevaddr__T_247_mask = 1'h1;
  assign mtlbptevaddr__T_247_en = ~io_rst_n;
  assign mtlbptevaddr__T_251_data = 32'h0;
  assign mtlbptevaddr__T_251_addr = 4'he;
  assign mtlbptevaddr__T_251_mask = 1'h1;
  assign mtlbptevaddr__T_251_en = ~io_rst_n;
  assign mtlbptevaddr__T_255_data = 32'h0;
  assign mtlbptevaddr__T_255_addr = 4'hf;
  assign mtlbptevaddr__T_255_mask = 1'h1;
  assign mtlbptevaddr__T_255_en = ~io_rst_n;
  assign mtlbptevaddr__T_475_data = io_data_i;
  assign mtlbptevaddr__T_475_addr = mtlbindex;
  assign mtlbptevaddr__T_475_mask = 1'h1;
  assign mtlbptevaddr__T_475_en = io_rst_n ? _GEN_1524 : 1'h0;
  assign _T_1 = mstatus_fs == 2'h3; // @[CSR.scala 76:53]
  assign _T_3 = io_prv_o < 2'h3; // @[CSR.scala 135:19]
  assign _T_4 = io_prv_o == 2'h3; // @[CSR.scala 135:47]
  assign _T_6 = _T_4 & mstatus_mie; // @[CSR.scala 135:63]
  assign _T_7 = _T_3 | _T_6; // @[CSR.scala 135:34]
  assign m_intr_globally_enabled = io_not_stall_i & _T_7; // @[CSR.scala 135:5]
  assign _T_9 = io_prv_o < 2'h1; // @[CSR.scala 140:19]
  assign _T_10 = io_prv_o == 2'h1; // @[CSR.scala 140:47]
  assign _T_12 = _T_10 & mstatus_sie; // @[CSR.scala 140:63]
  assign _T_13 = _T_9 | _T_12; // @[CSR.scala 140:34]
  assign s_intr_globally_enabled = io_not_stall_i & _T_13; // @[CSR.scala 140:5]
  assign _T_14 = mip_mtip & mie_mtie; // @[CSR.scala 144:31]
  assign _T_15 = _T_14 & m_intr_globally_enabled; // @[CSR.scala 144:42]
  assign m_mtime_intr = _T_15 & ~mideleg[7]; // @[CSR.scala 144:75]
  assign _T_18 = mip_msip & mie_msie; // @[CSR.scala 145:31]
  assign _T_19 = _T_18 & m_intr_globally_enabled; // @[CSR.scala 145:42]
  assign m_msoft_intr = _T_19 & ~mideleg[3]; // @[CSR.scala 145:75]
  assign _T_22 = mip_meip & mie_meie; // @[CSR.scala 146:31]
  assign _T_23 = _T_22 & m_intr_globally_enabled; // @[CSR.scala 146:42]
  assign m_mextr_intr = _T_23 & ~mideleg[11]; // @[CSR.scala 146:75]
  assign _T_26 = mip_stip & mie_stie; // @[CSR.scala 147:31]
  assign _T_27 = _T_26 & m_intr_globally_enabled; // @[CSR.scala 147:42]
  assign m_stime_intr = _T_27 & ~mideleg[5]; // @[CSR.scala 147:75]
  assign _T_30 = mip_ssip & mie_ssie; // @[CSR.scala 148:31]
  assign _T_31 = _T_30 & m_intr_globally_enabled; // @[CSR.scala 148:42]
  assign m_ssoft_intr = _T_31 & ~mideleg[1]; // @[CSR.scala 148:75]
  assign _T_34 = m_mtime_intr | m_msoft_intr; // @[CSR.scala 150:29]
  assign _T_35 = _T_34 | m_mextr_intr; // @[CSR.scala 150:44]
  assign _T_36 = _T_35 | m_stime_intr; // @[CSR.scala 150:59]
  assign m_intr = _T_36 | m_ssoft_intr; // @[CSR.scala 150:74]
  assign _T_38 = _T_14 & s_intr_globally_enabled; // @[CSR.scala 152:42]
  assign s_mtime_intr = _T_38 & mideleg[7]; // @[CSR.scala 152:75]
  assign _T_41 = _T_18 & s_intr_globally_enabled; // @[CSR.scala 153:42]
  assign s_msoft_intr = _T_41 & mideleg[3]; // @[CSR.scala 153:75]
  assign _T_44 = _T_22 & s_intr_globally_enabled; // @[CSR.scala 154:42]
  assign s_mextr_intr = _T_44 & mideleg[11]; // @[CSR.scala 154:75]
  assign _T_47 = _T_26 & s_intr_globally_enabled; // @[CSR.scala 155:42]
  assign s_stime_intr = _T_47 & mideleg[5]; // @[CSR.scala 155:75]
  assign _T_50 = _T_30 & s_intr_globally_enabled; // @[CSR.scala 156:42]
  assign s_ssoft_intr = _T_50 & mideleg[1]; // @[CSR.scala 156:75]
  assign _T_52 = s_mtime_intr | s_msoft_intr; // @[CSR.scala 158:29]
  assign _T_53 = _T_52 | s_mextr_intr; // @[CSR.scala 158:44]
  assign _T_54 = _T_53 | s_stime_intr; // @[CSR.scala 158:59]
  assign s_intr = _T_54 | s_ssoft_intr; // @[CSR.scala 158:74]
  assign _T_57 = io_not_stall_i & io_excepttype_i[0]; // @[CSR.scala 160:60]
  assign m_inst_misaligned_trap = _T_57 & ~medeleg[0]; // @[CSR.scala 160:110]
  assign _T_60 = {{1'd0}, io_excepttype_i[31:1]}; // @[CSR.scala 162:77]
  assign _T_62 = io_not_stall_i & _T_60[0]; // @[CSR.scala 162:60]
  assign m_inst_access_fault_trap = _T_62 & ~medeleg[1]; // @[CSR.scala 162:110]
  assign _T_65 = {{2'd0}, io_excepttype_i[31:2]}; // @[CSR.scala 164:77]
  assign _T_67 = io_not_stall_i & _T_65[0]; // @[CSR.scala 164:60]
  assign m_inst_illegal_trap = _T_67 & ~medeleg[2]; // @[CSR.scala 164:110]
  assign _T_70 = {{3'd0}, io_excepttype_i[31:3]}; // @[CSR.scala 166:77]
  assign _T_72 = io_not_stall_i & _T_70[0]; // @[CSR.scala 166:60]
  assign m_break_trap = _T_72 & ~medeleg[3]; // @[CSR.scala 166:110]
  assign _T_75 = {{4'd0}, io_excepttype_i[31:4]}; // @[CSR.scala 168:77]
  assign _T_77 = io_not_stall_i & _T_75[0]; // @[CSR.scala 168:60]
  assign m_load_misaligned_trap = _T_77 & ~medeleg[4]; // @[CSR.scala 168:110]
  assign _T_80 = {{5'd0}, io_excepttype_i[31:5]}; // @[CSR.scala 170:77]
  assign _T_82 = io_not_stall_i & _T_80[0]; // @[CSR.scala 170:60]
  assign m_load_access_fault_trap = _T_82 & ~medeleg[5]; // @[CSR.scala 170:110]
  assign _T_85 = {{6'd0}, io_excepttype_i[31:6]}; // @[CSR.scala 172:77]
  assign _T_87 = io_not_stall_i & _T_85[0]; // @[CSR.scala 172:60]
  assign m_store_misaligned_trap = _T_87 & ~medeleg[6]; // @[CSR.scala 172:110]
  assign _T_90 = {{7'd0}, io_excepttype_i[31:7]}; // @[CSR.scala 174:77]
  assign _T_92 = io_not_stall_i & _T_90[0]; // @[CSR.scala 174:60]
  assign m_store_access_fault_trap = _T_92 & ~medeleg[7]; // @[CSR.scala 174:110]
  assign _T_95 = {{8'd0}, io_excepttype_i[31:8]}; // @[CSR.scala 176:77]
  assign _T_97 = io_not_stall_i & _T_95[0]; // @[CSR.scala 176:60]
  assign m_ecall_from_u_trap = _T_97 & ~medeleg[8]; // @[CSR.scala 176:110]
  assign _T_100 = {{9'd0}, io_excepttype_i[31:9]}; // @[CSR.scala 178:77]
  assign _T_102 = io_not_stall_i & _T_100[0]; // @[CSR.scala 178:60]
  assign m_ecall_from_s_trap = _T_102 & ~medeleg[9]; // @[CSR.scala 178:110]
  assign _T_105 = {{11'd0}, io_excepttype_i[31:11]}; // @[CSR.scala 180:77]
  assign m_ecall_from_m_trap = io_not_stall_i & _T_105[0]; // @[CSR.scala 180:60]
  assign _T_107 = m_inst_misaligned_trap | m_inst_access_fault_trap; // @[CSR.scala 183:30]
  assign _T_108 = _T_107 | m_inst_illegal_trap; // @[CSR.scala 184:32]
  assign _T_109 = _T_108 | m_break_trap; // @[CSR.scala 185:27]
  assign _T_110 = _T_109 | m_load_misaligned_trap; // @[CSR.scala 186:20]
  assign _T_111 = _T_110 | m_load_access_fault_trap; // @[CSR.scala 187:30]
  assign _T_112 = _T_111 | m_store_misaligned_trap; // @[CSR.scala 188:32]
  assign _T_113 = _T_112 | m_store_access_fault_trap; // @[CSR.scala 189:31]
  assign _T_114 = _T_113 | m_ecall_from_u_trap; // @[CSR.scala 190:33]
  assign _T_115 = _T_114 | m_ecall_from_s_trap; // @[CSR.scala 191:27]
  assign m_trap = _T_115 | m_ecall_from_m_trap; // @[CSR.scala 192:27]
  assign _T_116 = {{15'd0}, io_excepttype_i[31:15]}; // @[CSR.scala 195:67]
  assign eret_from_m_trap = io_not_stall_i & _T_116[0]; // @[CSR.scala 195:50]
  assign _T_118 = {{13'd0}, io_excepttype_i[31:13]}; // @[CSR.scala 196:67]
  assign eret_from_s_trap = io_not_stall_i & _T_118[0]; // @[CSR.scala 196:50]
  assign _T_120 = {{21'd0}, io_excepttype_i[31:21]}; // @[CSR.scala 197:67]
  assign fence_i_trap = io_not_stall_i & _T_120[0]; // @[CSR.scala 197:50]
  assign s_inst_misaligned_trap = _T_57 & medeleg[0]; // @[CSR.scala 199:110]
  assign s_inst_access_fault_trap = _T_62 & medeleg[1]; // @[CSR.scala 201:110]
  assign s_inst_illegal_trap = _T_67 & medeleg[2]; // @[CSR.scala 203:110]
  assign s_break_trap = _T_72 & medeleg[3]; // @[CSR.scala 205:110]
  assign s_load_misaligned_trap = _T_77 & medeleg[4]; // @[CSR.scala 207:110]
  assign s_load_access_fault_trap = _T_82 & medeleg[5]; // @[CSR.scala 209:110]
  assign s_store_misaligned_trap = _T_87 & medeleg[6]; // @[CSR.scala 211:110]
  assign s_store_access_fault_trap = _T_92 & medeleg[7]; // @[CSR.scala 213:110]
  assign s_ecall_from_u_trap = _T_97 & medeleg[8]; // @[CSR.scala 215:110]
  assign s_ecall_from_s_trap = _T_102 & medeleg[9]; // @[CSR.scala 217:110]
  assign _T_162 = s_inst_misaligned_trap | s_inst_access_fault_trap; // @[CSR.scala 220:30]
  assign _T_163 = _T_162 | s_inst_illegal_trap; // @[CSR.scala 221:32]
  assign _T_164 = _T_163 | s_break_trap; // @[CSR.scala 222:27]
  assign _T_165 = _T_164 | s_load_misaligned_trap; // @[CSR.scala 223:20]
  assign _T_166 = _T_165 | s_load_access_fault_trap; // @[CSR.scala 224:30]
  assign _T_167 = _T_166 | s_store_misaligned_trap; // @[CSR.scala 225:32]
  assign _T_168 = _T_167 | s_store_access_fault_trap; // @[CSR.scala 226:31]
  assign _T_169 = _T_168 | s_ecall_from_u_trap; // @[CSR.scala 227:33]
  assign s_trap = _T_169 | s_ecall_from_s_trap; // @[CSR.scala 228:27]
  assign _T_172 = {mtvec_addr,1'h0}; // @[Cat.scala 29:58]
  assign _T_174 = {stvec_addr,1'h0}; // @[Cat.scala 29:58]
  assign _T_180 = {sepc_addr,1'h0}; // @[Cat.scala 29:58]
  assign _GEN_2048 = {{1'd0}, mstatus_spp}; // @[Conditional.scala 37:30]
  assign _T_181 = 2'h0 == _GEN_2048; // @[Conditional.scala 37:30]
  assign _T_182 = 2'h1 == _GEN_2048; // @[Conditional.scala 37:30]
  assign _T_184 = {mepc_addr,1'h0}; // @[Cat.scala 29:58]
  assign _T_185 = 2'h0 == mstatus_mpp; // @[Conditional.scala 37:30]
  assign _T_186 = 2'h1 == mstatus_mpp; // @[Conditional.scala 37:30]
  assign _T_187 = 2'h3 == mstatus_mpp; // @[Conditional.scala 37:30]
  assign _T_190 = io_current_inst_addr_i + 32'h4; // @[CSR.scala 277:55]
  assign _GEN_6 = fence_i_trap ? _T_190 : 32'h0; // @[CSR.scala 275:36]
  assign _GEN_7 = eret_from_m_trap | fence_i_trap; // @[CSR.scala 267:40]
  assign _GEN_8 = eret_from_m_trap ? {{1'd0}, _T_184} : _GEN_6; // @[CSR.scala 267:40]
  assign _GEN_10 = eret_from_s_trap | _GEN_7; // @[CSR.scala 260:40]
  assign _GEN_11 = eret_from_s_trap ? {{1'd0}, _T_180} : _GEN_8; // @[CSR.scala 260:40]
  assign _GEN_13 = s_trap | _GEN_10; // @[CSR.scala 256:30]
  assign _GEN_14 = s_trap ? {{1'd0}, _T_174} : _GEN_11; // @[CSR.scala 256:30]
  assign _GEN_16 = m_trap | _GEN_13; // @[CSR.scala 252:30]
  assign _GEN_17 = m_trap ? {{1'd0}, _T_172} : _GEN_14; // @[CSR.scala 252:30]
  assign _GEN_19 = s_intr | _GEN_16; // @[CSR.scala 248:30]
  assign _GEN_20 = s_intr ? {{1'd0}, _T_174} : _GEN_17; // @[CSR.scala 248:30]
  assign _GEN_22 = m_intr | _GEN_19; // @[CSR.scala 244:24]
  assign _GEN_23 = m_intr ? {{1'd0}, _T_172} : _GEN_20; // @[CSR.scala 244:24]
  assign _GEN_28 = m_mextr_intr | mcause_intr; // @[CSR.scala 365:37]
  assign _GEN_29 = m_mextr_intr ? 4'hb : mcause_code; // @[CSR.scala 365:37]
  assign _GEN_30 = m_mtime_intr | _GEN_28; // @[CSR.scala 362:37]
  assign _GEN_31 = m_mtime_intr ? 4'h7 : _GEN_29; // @[CSR.scala 362:37]
  assign _GEN_32 = m_stime_intr | _GEN_30; // @[CSR.scala 359:37]
  assign _GEN_33 = m_stime_intr ? 4'h5 : _GEN_31; // @[CSR.scala 359:37]
  assign _GEN_34 = m_msoft_intr | _GEN_32; // @[CSR.scala 356:37]
  assign _GEN_35 = m_msoft_intr ? 4'h3 : _GEN_33; // @[CSR.scala 356:37]
  assign _GEN_36 = m_ssoft_intr | _GEN_34; // @[CSR.scala 353:31]
  assign _GEN_37 = m_ssoft_intr ? 4'h1 : _GEN_35; // @[CSR.scala 353:31]
  assign _T_264 = 2'h0 == io_prv_o; // @[Conditional.scala 37:30]
  assign _T_265 = 2'h1 == io_prv_o; // @[Conditional.scala 37:30]
  assign _T_266 = 2'h3 == io_prv_o; // @[Conditional.scala 37:30]
  assign _GEN_44 = s_mextr_intr | scause_intr; // @[CSR.scala 399:37]
  assign _GEN_45 = s_mextr_intr ? 4'h5 : scause_code; // @[CSR.scala 399:37]
  assign _GEN_46 = s_mtime_intr | _GEN_44; // @[CSR.scala 396:37]
  assign _GEN_47 = s_mtime_intr ? 4'h5 : _GEN_45; // @[CSR.scala 396:37]
  assign _GEN_48 = s_stime_intr | _GEN_46; // @[CSR.scala 393:37]
  assign _GEN_49 = s_stime_intr ? 4'h5 : _GEN_47; // @[CSR.scala 393:37]
  assign _GEN_50 = s_msoft_intr | _GEN_48; // @[CSR.scala 390:37]
  assign _GEN_51 = s_msoft_intr ? 4'h1 : _GEN_49; // @[CSR.scala 390:37]
  assign _GEN_52 = s_ssoft_intr | _GEN_50; // @[CSR.scala 387:31]
  assign _GEN_53 = s_ssoft_intr ? 4'h1 : _GEN_51; // @[CSR.scala 387:31]
  assign _GEN_56 = _T_265 ? 2'h1 : {{1'd0}, mstatus_spp}; // @[Conditional.scala 39:67]
  assign _GEN_57 = _T_264 ? 2'h0 : _GEN_56; // @[Conditional.scala 40:58]
  assign _GEN_59 = m_ecall_from_m_trap ? 4'hb : mcause_code; // @[CSR.scala 455:44]
  assign _GEN_61 = m_ecall_from_s_trap ? 4'h9 : _GEN_59; // @[CSR.scala 452:44]
  assign _GEN_63 = m_ecall_from_u_trap ? 4'h8 : _GEN_61; // @[CSR.scala 449:44]
  assign _GEN_65 = m_store_access_fault_trap ? 4'h7 : _GEN_63; // @[CSR.scala 445:50]
  assign _GEN_68 = m_store_misaligned_trap ? 4'h6 : _GEN_65; // @[CSR.scala 441:48]
  assign _GEN_71 = m_load_access_fault_trap ? 4'h5 : _GEN_68; // @[CSR.scala 437:49]
  assign _GEN_74 = m_load_misaligned_trap ? 4'h4 : _GEN_71; // @[CSR.scala 433:47]
  assign _GEN_77 = m_break_trap ? 4'h3 : _GEN_74; // @[CSR.scala 430:37]
  assign _GEN_80 = m_inst_illegal_trap ? 4'h2 : _GEN_77; // @[CSR.scala 427:44]
  assign _GEN_83 = m_inst_access_fault_trap ? 4'h1 : _GEN_80; // @[CSR.scala 423:49]
  assign _GEN_86 = m_inst_misaligned_trap ? 4'h0 : _GEN_83; // @[CSR.scala 419:41]
  assign _GEN_95 = s_ecall_from_s_trap ? 4'h9 : mcause_code; // @[CSR.scala 510:44]
  assign _GEN_97 = s_ecall_from_u_trap ? 4'h8 : _GEN_95; // @[CSR.scala 507:44]
  assign _GEN_99 = s_store_access_fault_trap ? 4'h7 : _GEN_97; // @[CSR.scala 503:50]
  assign _GEN_102 = s_store_misaligned_trap ? 4'h6 : _GEN_99; // @[CSR.scala 499:48]
  assign _GEN_105 = s_load_access_fault_trap ? 4'h5 : _GEN_102; // @[CSR.scala 495:49]
  assign _GEN_108 = s_load_misaligned_trap ? 4'h4 : _GEN_105; // @[CSR.scala 491:47]
  assign _GEN_111 = s_break_trap ? 4'h3 : _GEN_108; // @[CSR.scala 488:37]
  assign _GEN_114 = s_inst_illegal_trap ? 4'h2 : _GEN_111; // @[CSR.scala 485:44]
  assign _GEN_117 = s_inst_access_fault_trap ? 4'h1 : _GEN_114; // @[CSR.scala 481:49]
  assign _GEN_120 = s_inst_misaligned_trap ? 4'h0 : _GEN_117; // @[CSR.scala 477:41]
  assign _GEN_127 = _T_182 | mstatus_spie; // @[Conditional.scala 39:67]
  assign _GEN_128 = _T_182 ? 1'h0 : mstatus_spp; // @[Conditional.scala 39:67]
  assign _GEN_129 = _T_181 | _GEN_127; // @[Conditional.scala 40:58]
  assign _GEN_130 = _T_181 ? 1'h0 : _GEN_128; // @[Conditional.scala 40:58]
  assign _GEN_133 = _T_187 | mstatus_mpie; // @[Conditional.scala 39:67]
  assign _GEN_136 = _T_186 | _GEN_133; // @[Conditional.scala 39:67]
  assign _GEN_138 = _T_185 | _GEN_136; // @[Conditional.scala 40:58]
  assign _T_325 = 12'h300 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_327 = 5'h0 == io_data_i[28:24]; // @[Conditional.scala 37:30]
  assign _T_328 = 5'h8 == io_data_i[28:24]; // @[Conditional.scala 37:30]
  assign _T_329 = _T_327 | _T_328; // @[Conditional.scala 37:55]
  assign _T_335 = 2'h3 == io_data_i[12:11]; // @[Conditional.scala 37:30]
  assign _T_336 = 2'h1 == io_data_i[12:11]; // @[Conditional.scala 37:30]
  assign _T_337 = 2'h0 == io_data_i[12:11]; // @[Conditional.scala 37:30]
  assign _T_338 = _T_335 | _T_336; // @[Conditional.scala 37:55]
  assign _T_339 = _T_338 | _T_337; // @[Conditional.scala 37:55]
  assign _T_342 = {1'h0,io_data_i[8]}; // @[Cat.scala 29:58]
  assign _T_343 = 2'h1 == _T_342; // @[Conditional.scala 37:30]
  assign _T_344 = 2'h0 == _T_342; // @[Conditional.scala 37:30]
  assign _T_345 = _T_343 | _T_344; // @[Conditional.scala 37:55]
  assign _GEN_143 = _T_345 ? io_data_i[8] : mstatus_spp; // @[Conditional.scala 40:58]
  assign _T_351 = 12'h344 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_354 = 12'h304 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_360 = 12'h321 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_362 = 12'h320 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_364 = 12'h340 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_365 = 12'h341 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_367 = 12'h305 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_369 = 12'h302 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_371 = 12'h303 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_373 = 12'h342 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_376 = {io_data_i[31],io_data_i[3:0]}; // @[Cat.scala 29:58]
  assign _T_377 = 5'h0 == _T_376; // @[Conditional.scala 37:30]
  assign _T_378 = 5'h1 == _T_376; // @[Conditional.scala 37:30]
  assign _T_379 = 5'h2 == _T_376; // @[Conditional.scala 37:30]
  assign _T_380 = 5'h3 == _T_376; // @[Conditional.scala 37:30]
  assign _T_381 = 5'h4 == _T_376; // @[Conditional.scala 37:30]
  assign _T_382 = 5'h5 == _T_376; // @[Conditional.scala 37:30]
  assign _T_383 = 5'h6 == _T_376; // @[Conditional.scala 37:30]
  assign _T_384 = 5'h7 == _T_376; // @[Conditional.scala 37:30]
  assign _T_385 = 5'h8 == _T_376; // @[Conditional.scala 37:30]
  assign _T_386 = 5'h9 == _T_376; // @[Conditional.scala 37:30]
  assign _T_387 = 5'ha == _T_376; // @[Conditional.scala 37:30]
  assign _T_388 = 5'hb == _T_376; // @[Conditional.scala 37:30]
  assign _T_389 = 5'h11 == _T_376; // @[Conditional.scala 37:30]
  assign _T_390 = 5'h13 == _T_376; // @[Conditional.scala 37:30]
  assign _T_391 = 5'h15 == _T_376; // @[Conditional.scala 37:30]
  assign _T_392 = 5'h17 == _T_376; // @[Conditional.scala 37:30]
  assign _T_393 = 5'h1b == _T_376; // @[Conditional.scala 37:30]
  assign _T_394 = _T_377 | _T_378; // @[Conditional.scala 37:55]
  assign _T_395 = _T_394 | _T_379; // @[Conditional.scala 37:55]
  assign _T_396 = _T_395 | _T_380; // @[Conditional.scala 37:55]
  assign _T_397 = _T_396 | _T_381; // @[Conditional.scala 37:55]
  assign _T_398 = _T_397 | _T_382; // @[Conditional.scala 37:55]
  assign _T_399 = _T_398 | _T_383; // @[Conditional.scala 37:55]
  assign _T_400 = _T_399 | _T_384; // @[Conditional.scala 37:55]
  assign _T_401 = _T_400 | _T_385; // @[Conditional.scala 37:55]
  assign _T_402 = _T_401 | _T_386; // @[Conditional.scala 37:55]
  assign _T_403 = _T_402 | _T_387; // @[Conditional.scala 37:55]
  assign _T_404 = _T_403 | _T_388; // @[Conditional.scala 37:55]
  assign _T_405 = _T_404 | _T_389; // @[Conditional.scala 37:55]
  assign _T_406 = _T_405 | _T_390; // @[Conditional.scala 37:55]
  assign _T_407 = _T_406 | _T_391; // @[Conditional.scala 37:55]
  assign _T_408 = _T_407 | _T_392; // @[Conditional.scala 37:55]
  assign _T_409 = _T_408 | _T_393; // @[Conditional.scala 37:55]
  assign _GEN_145 = _T_409 ? io_data_i[3:0] : mcause_code; // @[Conditional.scala 40:58]
  assign _T_412 = 12'h343 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_413 = 12'h100 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_423 = 12'h105 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_425 = 12'h144 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_428 = 12'h104 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_431 = 12'h140 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_432 = 12'h141 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_434 = 12'h142 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_459 = _T_402 | _T_389; // @[Conditional.scala 37:55]
  assign _T_460 = _T_459 | _T_391; // @[Conditional.scala 37:55]
  assign _GEN_148 = _T_460 ? io_data_i[3:0] : scause_code; // @[Conditional.scala 40:58]
  assign _T_463 = 12'h143 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_464 = 12'h180 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_466 = 12'h7c0 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_468 = 12'h7c1 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_470 = 12'h7c2 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_472 = 12'h7c3 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _T_474 = 12'h7c4 == io_waddr_i; // @[Conditional.scala 37:30]
  assign _GEN_161 = _T_472 ? 1'h0 : _T_474; // @[Conditional.scala 39:67]
  assign _GEN_171 = _T_470 ? 1'h0 : _T_472; // @[Conditional.scala 39:67]
  assign _GEN_176 = _T_470 ? 1'h0 : _GEN_161; // @[Conditional.scala 39:67]
  assign _GEN_186 = _T_468 ? 1'h0 : _T_470; // @[Conditional.scala 39:67]
  assign _GEN_191 = _T_468 ? 1'h0 : _GEN_171; // @[Conditional.scala 39:67]
  assign _GEN_196 = _T_468 ? 1'h0 : _GEN_176; // @[Conditional.scala 39:67]
  assign _GEN_199 = _T_466 ? io_data_i[3:0] : mtlbindex; // @[Conditional.scala 39:67]
  assign _GEN_200 = _T_466 ? 1'h0 : mtlbindex_update; // @[Conditional.scala 39:67]
  assign _GEN_203 = _T_466 ? 1'h0 : _T_468; // @[Conditional.scala 39:67]
  assign _GEN_208 = _T_466 ? 1'h0 : _GEN_186; // @[Conditional.scala 39:67]
  assign _GEN_213 = _T_466 ? 1'h0 : _GEN_191; // @[Conditional.scala 39:67]
  assign _GEN_218 = _T_466 ? 1'h0 : _GEN_196; // @[Conditional.scala 39:67]
  assign _GEN_221 = _T_464 ? io_data_i[21:0] : sptbr_ppn; // @[Conditional.scala 39:67]
  assign _GEN_222 = _T_464 ? mtlbindex : _GEN_199; // @[Conditional.scala 39:67]
  assign _GEN_223 = _T_464 ? mtlbindex_update : _GEN_200; // @[Conditional.scala 39:67]
  assign _GEN_226 = _T_464 ? 1'h0 : _GEN_203; // @[Conditional.scala 39:67]
  assign _GEN_231 = _T_464 ? 1'h0 : _GEN_208; // @[Conditional.scala 39:67]
  assign _GEN_236 = _T_464 ? 1'h0 : _GEN_213; // @[Conditional.scala 39:67]
  assign _GEN_241 = _T_464 ? 1'h0 : _GEN_218; // @[Conditional.scala 39:67]
  assign _GEN_245 = _T_463 ? sptbr_ppn : _GEN_221; // @[Conditional.scala 39:67]
  assign _GEN_246 = _T_463 ? mtlbindex : _GEN_222; // @[Conditional.scala 39:67]
  assign _GEN_247 = _T_463 ? mtlbindex_update : _GEN_223; // @[Conditional.scala 39:67]
  assign _GEN_250 = _T_463 ? 1'h0 : _GEN_226; // @[Conditional.scala 39:67]
  assign _GEN_255 = _T_463 ? 1'h0 : _GEN_231; // @[Conditional.scala 39:67]
  assign _GEN_260 = _T_463 ? 1'h0 : _GEN_236; // @[Conditional.scala 39:67]
  assign _GEN_265 = _T_463 ? 1'h0 : _GEN_241; // @[Conditional.scala 39:67]
  assign _GEN_269 = _T_434 ? _GEN_148 : scause_code; // @[Conditional.scala 39:67]
  assign _GEN_271 = _T_434 ? sptbr_ppn : _GEN_245; // @[Conditional.scala 39:67]
  assign _GEN_272 = _T_434 ? mtlbindex : _GEN_246; // @[Conditional.scala 39:67]
  assign _GEN_273 = _T_434 ? mtlbindex_update : _GEN_247; // @[Conditional.scala 39:67]
  assign _GEN_276 = _T_434 ? 1'h0 : _GEN_250; // @[Conditional.scala 39:67]
  assign _GEN_281 = _T_434 ? 1'h0 : _GEN_255; // @[Conditional.scala 39:67]
  assign _GEN_286 = _T_434 ? 1'h0 : _GEN_260; // @[Conditional.scala 39:67]
  assign _GEN_291 = _T_434 ? 1'h0 : _GEN_265; // @[Conditional.scala 39:67]
  assign _GEN_294 = _T_432 ? io_data_i[31:2] : sepc_addr; // @[Conditional.scala 39:67]
  assign _GEN_296 = _T_432 ? scause_code : _GEN_269; // @[Conditional.scala 39:67]
  assign _GEN_298 = _T_432 ? sptbr_ppn : _GEN_271; // @[Conditional.scala 39:67]
  assign _GEN_299 = _T_432 ? mtlbindex : _GEN_272; // @[Conditional.scala 39:67]
  assign _GEN_300 = _T_432 ? mtlbindex_update : _GEN_273; // @[Conditional.scala 39:67]
  assign _GEN_303 = _T_432 ? 1'h0 : _GEN_276; // @[Conditional.scala 39:67]
  assign _GEN_308 = _T_432 ? 1'h0 : _GEN_281; // @[Conditional.scala 39:67]
  assign _GEN_313 = _T_432 ? 1'h0 : _GEN_286; // @[Conditional.scala 39:67]
  assign _GEN_318 = _T_432 ? 1'h0 : _GEN_291; // @[Conditional.scala 39:67]
  assign _GEN_322 = _T_431 ? sepc_addr : _GEN_294; // @[Conditional.scala 39:67]
  assign _GEN_324 = _T_431 ? scause_code : _GEN_296; // @[Conditional.scala 39:67]
  assign _GEN_326 = _T_431 ? sptbr_ppn : _GEN_298; // @[Conditional.scala 39:67]
  assign _GEN_327 = _T_431 ? mtlbindex : _GEN_299; // @[Conditional.scala 39:67]
  assign _GEN_328 = _T_431 ? mtlbindex_update : _GEN_300; // @[Conditional.scala 39:67]
  assign _GEN_331 = _T_431 ? 1'h0 : _GEN_303; // @[Conditional.scala 39:67]
  assign _GEN_336 = _T_431 ? 1'h0 : _GEN_308; // @[Conditional.scala 39:67]
  assign _GEN_341 = _T_431 ? 1'h0 : _GEN_313; // @[Conditional.scala 39:67]
  assign _GEN_346 = _T_431 ? 1'h0 : _GEN_318; // @[Conditional.scala 39:67]
  assign _GEN_352 = _T_428 ? sepc_addr : _GEN_322; // @[Conditional.scala 39:67]
  assign _GEN_354 = _T_428 ? scause_code : _GEN_324; // @[Conditional.scala 39:67]
  assign _GEN_356 = _T_428 ? sptbr_ppn : _GEN_326; // @[Conditional.scala 39:67]
  assign _GEN_357 = _T_428 ? mtlbindex : _GEN_327; // @[Conditional.scala 39:67]
  assign _GEN_358 = _T_428 ? mtlbindex_update : _GEN_328; // @[Conditional.scala 39:67]
  assign _GEN_361 = _T_428 ? 1'h0 : _GEN_331; // @[Conditional.scala 39:67]
  assign _GEN_366 = _T_428 ? 1'h0 : _GEN_336; // @[Conditional.scala 39:67]
  assign _GEN_371 = _T_428 ? 1'h0 : _GEN_341; // @[Conditional.scala 39:67]
  assign _GEN_376 = _T_428 ? 1'h0 : _GEN_346; // @[Conditional.scala 39:67]
  assign _GEN_384 = _T_425 ? sepc_addr : _GEN_352; // @[Conditional.scala 39:67]
  assign _GEN_386 = _T_425 ? scause_code : _GEN_354; // @[Conditional.scala 39:67]
  assign _GEN_388 = _T_425 ? sptbr_ppn : _GEN_356; // @[Conditional.scala 39:67]
  assign _GEN_389 = _T_425 ? mtlbindex : _GEN_357; // @[Conditional.scala 39:67]
  assign _GEN_390 = _T_425 ? mtlbindex_update : _GEN_358; // @[Conditional.scala 39:67]
  assign _GEN_393 = _T_425 ? 1'h0 : _GEN_361; // @[Conditional.scala 39:67]
  assign _GEN_398 = _T_425 ? 1'h0 : _GEN_366; // @[Conditional.scala 39:67]
  assign _GEN_403 = _T_425 ? 1'h0 : _GEN_371; // @[Conditional.scala 39:67]
  assign _GEN_408 = _T_425 ? 1'h0 : _GEN_376; // @[Conditional.scala 39:67]
  assign _GEN_411 = _T_423 ? io_data_i[31:2] : stvec_addr; // @[Conditional.scala 39:67]
  assign _GEN_417 = _T_423 ? sepc_addr : _GEN_384; // @[Conditional.scala 39:67]
  assign _GEN_419 = _T_423 ? scause_code : _GEN_386; // @[Conditional.scala 39:67]
  assign _GEN_421 = _T_423 ? sptbr_ppn : _GEN_388; // @[Conditional.scala 39:67]
  assign _GEN_422 = _T_423 ? mtlbindex : _GEN_389; // @[Conditional.scala 39:67]
  assign _GEN_423 = _T_423 ? mtlbindex_update : _GEN_390; // @[Conditional.scala 39:67]
  assign _GEN_426 = _T_423 ? 1'h0 : _GEN_393; // @[Conditional.scala 39:67]
  assign _GEN_431 = _T_423 ? 1'h0 : _GEN_398; // @[Conditional.scala 39:67]
  assign _GEN_436 = _T_423 ? 1'h0 : _GEN_403; // @[Conditional.scala 39:67]
  assign _GEN_441 = _T_423 ? 1'h0 : _GEN_408; // @[Conditional.scala 39:67]
  assign _GEN_445 = _T_413 ? _GEN_143 : mstatus_spp; // @[Conditional.scala 39:67]
  assign _GEN_448 = _T_413 ? stvec_addr : _GEN_411; // @[Conditional.scala 39:67]
  assign _GEN_454 = _T_413 ? sepc_addr : _GEN_417; // @[Conditional.scala 39:67]
  assign _GEN_456 = _T_413 ? scause_code : _GEN_419; // @[Conditional.scala 39:67]
  assign _GEN_458 = _T_413 ? sptbr_ppn : _GEN_421; // @[Conditional.scala 39:67]
  assign _GEN_459 = _T_413 ? mtlbindex : _GEN_422; // @[Conditional.scala 39:67]
  assign _GEN_460 = _T_413 ? mtlbindex_update : _GEN_423; // @[Conditional.scala 39:67]
  assign _GEN_463 = _T_413 ? 1'h0 : _GEN_426; // @[Conditional.scala 39:67]
  assign _GEN_468 = _T_413 ? 1'h0 : _GEN_431; // @[Conditional.scala 39:67]
  assign _GEN_473 = _T_413 ? 1'h0 : _GEN_436; // @[Conditional.scala 39:67]
  assign _GEN_478 = _T_413 ? 1'h0 : _GEN_441; // @[Conditional.scala 39:67]
  assign _GEN_483 = _T_412 ? mstatus_spp : _GEN_445; // @[Conditional.scala 39:67]
  assign _GEN_486 = _T_412 ? stvec_addr : _GEN_448; // @[Conditional.scala 39:67]
  assign _GEN_492 = _T_412 ? sepc_addr : _GEN_454; // @[Conditional.scala 39:67]
  assign _GEN_494 = _T_412 ? scause_code : _GEN_456; // @[Conditional.scala 39:67]
  assign _GEN_496 = _T_412 ? sptbr_ppn : _GEN_458; // @[Conditional.scala 39:67]
  assign _GEN_497 = _T_412 ? mtlbindex : _GEN_459; // @[Conditional.scala 39:67]
  assign _GEN_498 = _T_412 ? mtlbindex_update : _GEN_460; // @[Conditional.scala 39:67]
  assign _GEN_501 = _T_412 ? 1'h0 : _GEN_463; // @[Conditional.scala 39:67]
  assign _GEN_506 = _T_412 ? 1'h0 : _GEN_468; // @[Conditional.scala 39:67]
  assign _GEN_511 = _T_412 ? 1'h0 : _GEN_473; // @[Conditional.scala 39:67]
  assign _GEN_516 = _T_412 ? 1'h0 : _GEN_478; // @[Conditional.scala 39:67]
  assign _GEN_520 = _T_373 ? _GEN_145 : mcause_code; // @[Conditional.scala 39:67]
  assign _GEN_523 = _T_373 ? mstatus_spp : _GEN_483; // @[Conditional.scala 39:67]
  assign _GEN_526 = _T_373 ? stvec_addr : _GEN_486; // @[Conditional.scala 39:67]
  assign _GEN_532 = _T_373 ? sepc_addr : _GEN_492; // @[Conditional.scala 39:67]
  assign _GEN_534 = _T_373 ? scause_code : _GEN_494; // @[Conditional.scala 39:67]
  assign _GEN_536 = _T_373 ? sptbr_ppn : _GEN_496; // @[Conditional.scala 39:67]
  assign _GEN_537 = _T_373 ? mtlbindex : _GEN_497; // @[Conditional.scala 39:67]
  assign _GEN_538 = _T_373 ? mtlbindex_update : _GEN_498; // @[Conditional.scala 39:67]
  assign _GEN_541 = _T_373 ? 1'h0 : _GEN_501; // @[Conditional.scala 39:67]
  assign _GEN_546 = _T_373 ? 1'h0 : _GEN_506; // @[Conditional.scala 39:67]
  assign _GEN_551 = _T_373 ? 1'h0 : _GEN_511; // @[Conditional.scala 39:67]
  assign _GEN_556 = _T_373 ? 1'h0 : _GEN_516; // @[Conditional.scala 39:67]
  assign _GEN_559 = _T_371 ? io_data_i[11:0] : mideleg; // @[Conditional.scala 39:67]
  assign _GEN_561 = _T_371 ? mcause_code : _GEN_520; // @[Conditional.scala 39:67]
  assign _GEN_564 = _T_371 ? mstatus_spp : _GEN_523; // @[Conditional.scala 39:67]
  assign _GEN_567 = _T_371 ? stvec_addr : _GEN_526; // @[Conditional.scala 39:67]
  assign _GEN_573 = _T_371 ? sepc_addr : _GEN_532; // @[Conditional.scala 39:67]
  assign _GEN_575 = _T_371 ? scause_code : _GEN_534; // @[Conditional.scala 39:67]
  assign _GEN_577 = _T_371 ? sptbr_ppn : _GEN_536; // @[Conditional.scala 39:67]
  assign _GEN_578 = _T_371 ? mtlbindex : _GEN_537; // @[Conditional.scala 39:67]
  assign _GEN_579 = _T_371 ? mtlbindex_update : _GEN_538; // @[Conditional.scala 39:67]
  assign _GEN_582 = _T_371 ? 1'h0 : _GEN_541; // @[Conditional.scala 39:67]
  assign _GEN_587 = _T_371 ? 1'h0 : _GEN_546; // @[Conditional.scala 39:67]
  assign _GEN_592 = _T_371 ? 1'h0 : _GEN_551; // @[Conditional.scala 39:67]
  assign _GEN_597 = _T_371 ? 1'h0 : _GEN_556; // @[Conditional.scala 39:67]
  assign _GEN_600 = _T_369 ? io_data_i[11:0] : medeleg; // @[Conditional.scala 39:67]
  assign _GEN_601 = _T_369 ? mideleg : _GEN_559; // @[Conditional.scala 39:67]
  assign _GEN_603 = _T_369 ? mcause_code : _GEN_561; // @[Conditional.scala 39:67]
  assign _GEN_606 = _T_369 ? mstatus_spp : _GEN_564; // @[Conditional.scala 39:67]
  assign _GEN_609 = _T_369 ? stvec_addr : _GEN_567; // @[Conditional.scala 39:67]
  assign _GEN_615 = _T_369 ? sepc_addr : _GEN_573; // @[Conditional.scala 39:67]
  assign _GEN_617 = _T_369 ? scause_code : _GEN_575; // @[Conditional.scala 39:67]
  assign _GEN_619 = _T_369 ? sptbr_ppn : _GEN_577; // @[Conditional.scala 39:67]
  assign _GEN_620 = _T_369 ? mtlbindex : _GEN_578; // @[Conditional.scala 39:67]
  assign _GEN_621 = _T_369 ? mtlbindex_update : _GEN_579; // @[Conditional.scala 39:67]
  assign _GEN_624 = _T_369 ? 1'h0 : _GEN_582; // @[Conditional.scala 39:67]
  assign _GEN_629 = _T_369 ? 1'h0 : _GEN_587; // @[Conditional.scala 39:67]
  assign _GEN_634 = _T_369 ? 1'h0 : _GEN_592; // @[Conditional.scala 39:67]
  assign _GEN_639 = _T_369 ? 1'h0 : _GEN_597; // @[Conditional.scala 39:67]
  assign _GEN_642 = _T_367 ? io_data_i[31:2] : mtvec_addr; // @[Conditional.scala 39:67]
  assign _GEN_643 = _T_367 ? medeleg : _GEN_600; // @[Conditional.scala 39:67]
  assign _GEN_644 = _T_367 ? mideleg : _GEN_601; // @[Conditional.scala 39:67]
  assign _GEN_646 = _T_367 ? mcause_code : _GEN_603; // @[Conditional.scala 39:67]
  assign _GEN_649 = _T_367 ? mstatus_spp : _GEN_606; // @[Conditional.scala 39:67]
  assign _GEN_652 = _T_367 ? stvec_addr : _GEN_609; // @[Conditional.scala 39:67]
  assign _GEN_658 = _T_367 ? sepc_addr : _GEN_615; // @[Conditional.scala 39:67]
  assign _GEN_660 = _T_367 ? scause_code : _GEN_617; // @[Conditional.scala 39:67]
  assign _GEN_662 = _T_367 ? sptbr_ppn : _GEN_619; // @[Conditional.scala 39:67]
  assign _GEN_663 = _T_367 ? mtlbindex : _GEN_620; // @[Conditional.scala 39:67]
  assign _GEN_664 = _T_367 ? mtlbindex_update : _GEN_621; // @[Conditional.scala 39:67]
  assign _GEN_667 = _T_367 ? 1'h0 : _GEN_624; // @[Conditional.scala 39:67]
  assign _GEN_672 = _T_367 ? 1'h0 : _GEN_629; // @[Conditional.scala 39:67]
  assign _GEN_677 = _T_367 ? 1'h0 : _GEN_634; // @[Conditional.scala 39:67]
  assign _GEN_682 = _T_367 ? 1'h0 : _GEN_639; // @[Conditional.scala 39:67]
  assign _GEN_685 = _T_365 ? io_data_i[31:2] : mepc_addr; // @[Conditional.scala 39:67]
  assign _GEN_686 = _T_365 ? mtvec_addr : _GEN_642; // @[Conditional.scala 39:67]
  assign _GEN_687 = _T_365 ? medeleg : _GEN_643; // @[Conditional.scala 39:67]
  assign _GEN_688 = _T_365 ? mideleg : _GEN_644; // @[Conditional.scala 39:67]
  assign _GEN_690 = _T_365 ? mcause_code : _GEN_646; // @[Conditional.scala 39:67]
  assign _GEN_693 = _T_365 ? mstatus_spp : _GEN_649; // @[Conditional.scala 39:67]
  assign _GEN_696 = _T_365 ? stvec_addr : _GEN_652; // @[Conditional.scala 39:67]
  assign _GEN_702 = _T_365 ? sepc_addr : _GEN_658; // @[Conditional.scala 39:67]
  assign _GEN_704 = _T_365 ? scause_code : _GEN_660; // @[Conditional.scala 39:67]
  assign _GEN_706 = _T_365 ? sptbr_ppn : _GEN_662; // @[Conditional.scala 39:67]
  assign _GEN_707 = _T_365 ? mtlbindex : _GEN_663; // @[Conditional.scala 39:67]
  assign _GEN_708 = _T_365 ? mtlbindex_update : _GEN_664; // @[Conditional.scala 39:67]
  assign _GEN_711 = _T_365 ? 1'h0 : _GEN_667; // @[Conditional.scala 39:67]
  assign _GEN_716 = _T_365 ? 1'h0 : _GEN_672; // @[Conditional.scala 39:67]
  assign _GEN_721 = _T_365 ? 1'h0 : _GEN_677; // @[Conditional.scala 39:67]
  assign _GEN_726 = _T_365 ? 1'h0 : _GEN_682; // @[Conditional.scala 39:67]
  assign _GEN_730 = _T_364 ? mepc_addr : _GEN_685; // @[Conditional.scala 39:67]
  assign _GEN_731 = _T_364 ? mtvec_addr : _GEN_686; // @[Conditional.scala 39:67]
  assign _GEN_732 = _T_364 ? medeleg : _GEN_687; // @[Conditional.scala 39:67]
  assign _GEN_733 = _T_364 ? mideleg : _GEN_688; // @[Conditional.scala 39:67]
  assign _GEN_735 = _T_364 ? mcause_code : _GEN_690; // @[Conditional.scala 39:67]
  assign _GEN_738 = _T_364 ? mstatus_spp : _GEN_693; // @[Conditional.scala 39:67]
  assign _GEN_741 = _T_364 ? stvec_addr : _GEN_696; // @[Conditional.scala 39:67]
  assign _GEN_747 = _T_364 ? sepc_addr : _GEN_702; // @[Conditional.scala 39:67]
  assign _GEN_749 = _T_364 ? scause_code : _GEN_704; // @[Conditional.scala 39:67]
  assign _GEN_751 = _T_364 ? sptbr_ppn : _GEN_706; // @[Conditional.scala 39:67]
  assign _GEN_752 = _T_364 ? mtlbindex : _GEN_707; // @[Conditional.scala 39:67]
  assign _GEN_753 = _T_364 ? mtlbindex_update : _GEN_708; // @[Conditional.scala 39:67]
  assign _GEN_756 = _T_364 ? 1'h0 : _GEN_711; // @[Conditional.scala 39:67]
  assign _GEN_761 = _T_364 ? 1'h0 : _GEN_716; // @[Conditional.scala 39:67]
  assign _GEN_766 = _T_364 ? 1'h0 : _GEN_721; // @[Conditional.scala 39:67]
  assign _GEN_771 = _T_364 ? 1'h0 : _GEN_726; // @[Conditional.scala 39:67]
  assign _GEN_776 = _T_362 ? mepc_addr : _GEN_730; // @[Conditional.scala 39:67]
  assign _GEN_777 = _T_362 ? mtvec_addr : _GEN_731; // @[Conditional.scala 39:67]
  assign _GEN_778 = _T_362 ? medeleg : _GEN_732; // @[Conditional.scala 39:67]
  assign _GEN_779 = _T_362 ? mideleg : _GEN_733; // @[Conditional.scala 39:67]
  assign _GEN_781 = _T_362 ? mcause_code : _GEN_735; // @[Conditional.scala 39:67]
  assign _GEN_784 = _T_362 ? mstatus_spp : _GEN_738; // @[Conditional.scala 39:67]
  assign _GEN_787 = _T_362 ? stvec_addr : _GEN_741; // @[Conditional.scala 39:67]
  assign _GEN_793 = _T_362 ? sepc_addr : _GEN_747; // @[Conditional.scala 39:67]
  assign _GEN_795 = _T_362 ? scause_code : _GEN_749; // @[Conditional.scala 39:67]
  assign _GEN_797 = _T_362 ? sptbr_ppn : _GEN_751; // @[Conditional.scala 39:67]
  assign _GEN_798 = _T_362 ? mtlbindex : _GEN_752; // @[Conditional.scala 39:67]
  assign _GEN_799 = _T_362 ? mtlbindex_update : _GEN_753; // @[Conditional.scala 39:67]
  assign _GEN_802 = _T_362 ? 1'h0 : _GEN_756; // @[Conditional.scala 39:67]
  assign _GEN_807 = _T_362 ? 1'h0 : _GEN_761; // @[Conditional.scala 39:67]
  assign _GEN_812 = _T_362 ? 1'h0 : _GEN_766; // @[Conditional.scala 39:67]
  assign _GEN_817 = _T_362 ? 1'h0 : _GEN_771; // @[Conditional.scala 39:67]
  assign _GEN_823 = _T_360 ? mepc_addr : _GEN_776; // @[Conditional.scala 39:67]
  assign _GEN_824 = _T_360 ? mtvec_addr : _GEN_777; // @[Conditional.scala 39:67]
  assign _GEN_825 = _T_360 ? medeleg : _GEN_778; // @[Conditional.scala 39:67]
  assign _GEN_826 = _T_360 ? mideleg : _GEN_779; // @[Conditional.scala 39:67]
  assign _GEN_828 = _T_360 ? mcause_code : _GEN_781; // @[Conditional.scala 39:67]
  assign _GEN_831 = _T_360 ? mstatus_spp : _GEN_784; // @[Conditional.scala 39:67]
  assign _GEN_834 = _T_360 ? stvec_addr : _GEN_787; // @[Conditional.scala 39:67]
  assign _GEN_840 = _T_360 ? sepc_addr : _GEN_793; // @[Conditional.scala 39:67]
  assign _GEN_842 = _T_360 ? scause_code : _GEN_795; // @[Conditional.scala 39:67]
  assign _GEN_844 = _T_360 ? sptbr_ppn : _GEN_797; // @[Conditional.scala 39:67]
  assign _GEN_845 = _T_360 ? mtlbindex : _GEN_798; // @[Conditional.scala 39:67]
  assign _GEN_846 = _T_360 ? mtlbindex_update : _GEN_799; // @[Conditional.scala 39:67]
  assign _GEN_849 = _T_360 ? 1'h0 : _GEN_802; // @[Conditional.scala 39:67]
  assign _GEN_854 = _T_360 ? 1'h0 : _GEN_807; // @[Conditional.scala 39:67]
  assign _GEN_859 = _T_360 ? 1'h0 : _GEN_812; // @[Conditional.scala 39:67]
  assign _GEN_864 = _T_360 ? 1'h0 : _GEN_817; // @[Conditional.scala 39:67]
  assign _GEN_875 = _T_354 ? mepc_addr : _GEN_823; // @[Conditional.scala 39:67]
  assign _GEN_876 = _T_354 ? mtvec_addr : _GEN_824; // @[Conditional.scala 39:67]
  assign _GEN_877 = _T_354 ? medeleg : _GEN_825; // @[Conditional.scala 39:67]
  assign _GEN_878 = _T_354 ? mideleg : _GEN_826; // @[Conditional.scala 39:67]
  assign _GEN_880 = _T_354 ? mcause_code : _GEN_828; // @[Conditional.scala 39:67]
  assign _GEN_883 = _T_354 ? mstatus_spp : _GEN_831; // @[Conditional.scala 39:67]
  assign _GEN_886 = _T_354 ? stvec_addr : _GEN_834; // @[Conditional.scala 39:67]
  assign _GEN_890 = _T_354 ? sepc_addr : _GEN_840; // @[Conditional.scala 39:67]
  assign _GEN_892 = _T_354 ? scause_code : _GEN_842; // @[Conditional.scala 39:67]
  assign _GEN_894 = _T_354 ? sptbr_ppn : _GEN_844; // @[Conditional.scala 39:67]
  assign _GEN_895 = _T_354 ? mtlbindex : _GEN_845; // @[Conditional.scala 39:67]
  assign _GEN_896 = _T_354 ? mtlbindex_update : _GEN_846; // @[Conditional.scala 39:67]
  assign _GEN_899 = _T_354 ? 1'h0 : _GEN_849; // @[Conditional.scala 39:67]
  assign _GEN_904 = _T_354 ? 1'h0 : _GEN_854; // @[Conditional.scala 39:67]
  assign _GEN_909 = _T_354 ? 1'h0 : _GEN_859; // @[Conditional.scala 39:67]
  assign _GEN_914 = _T_354 ? 1'h0 : _GEN_864; // @[Conditional.scala 39:67]
  assign _GEN_927 = _T_351 ? mepc_addr : _GEN_875; // @[Conditional.scala 39:67]
  assign _GEN_928 = _T_351 ? mtvec_addr : _GEN_876; // @[Conditional.scala 39:67]
  assign _GEN_929 = _T_351 ? medeleg : _GEN_877; // @[Conditional.scala 39:67]
  assign _GEN_930 = _T_351 ? mideleg : _GEN_878; // @[Conditional.scala 39:67]
  assign _GEN_932 = _T_351 ? mcause_code : _GEN_880; // @[Conditional.scala 39:67]
  assign _GEN_935 = _T_351 ? mstatus_spp : _GEN_883; // @[Conditional.scala 39:67]
  assign _GEN_938 = _T_351 ? stvec_addr : _GEN_886; // @[Conditional.scala 39:67]
  assign _GEN_940 = _T_351 ? sepc_addr : _GEN_890; // @[Conditional.scala 39:67]
  assign _GEN_942 = _T_351 ? scause_code : _GEN_892; // @[Conditional.scala 39:67]
  assign _GEN_944 = _T_351 ? sptbr_ppn : _GEN_894; // @[Conditional.scala 39:67]
  assign _GEN_945 = _T_351 ? mtlbindex : _GEN_895; // @[Conditional.scala 39:67]
  assign _GEN_946 = _T_351 ? mtlbindex_update : _GEN_896; // @[Conditional.scala 39:67]
  assign _GEN_949 = _T_351 ? 1'h0 : _GEN_899; // @[Conditional.scala 39:67]
  assign _GEN_954 = _T_351 ? 1'h0 : _GEN_904; // @[Conditional.scala 39:67]
  assign _GEN_959 = _T_351 ? 1'h0 : _GEN_909; // @[Conditional.scala 39:67]
  assign _GEN_964 = _T_351 ? 1'h0 : _GEN_914; // @[Conditional.scala 39:67]
  assign _GEN_972 = _T_325 ? _GEN_143 : _GEN_935; // @[Conditional.scala 40:58]
  assign _GEN_987 = _T_325 ? mepc_addr : _GEN_927; // @[Conditional.scala 40:58]
  assign _GEN_988 = _T_325 ? mtvec_addr : _GEN_928; // @[Conditional.scala 40:58]
  assign _GEN_989 = _T_325 ? medeleg : _GEN_929; // @[Conditional.scala 40:58]
  assign _GEN_990 = _T_325 ? mideleg : _GEN_930; // @[Conditional.scala 40:58]
  assign _GEN_992 = _T_325 ? mcause_code : _GEN_932; // @[Conditional.scala 40:58]
  assign _GEN_994 = _T_325 ? stvec_addr : _GEN_938; // @[Conditional.scala 40:58]
  assign _GEN_996 = _T_325 ? sepc_addr : _GEN_940; // @[Conditional.scala 40:58]
  assign _GEN_998 = _T_325 ? scause_code : _GEN_942; // @[Conditional.scala 40:58]
  assign _GEN_1000 = _T_325 ? sptbr_ppn : _GEN_944; // @[Conditional.scala 40:58]
  assign _GEN_1001 = _T_325 ? mtlbindex : _GEN_945; // @[Conditional.scala 40:58]
  assign _GEN_1002 = _T_325 ? mtlbindex_update : _GEN_946; // @[Conditional.scala 40:58]
  assign _GEN_1005 = _T_325 ? 1'h0 : _GEN_949; // @[Conditional.scala 40:58]
  assign _GEN_1010 = _T_325 ? 1'h0 : _GEN_954; // @[Conditional.scala 40:58]
  assign _GEN_1015 = _T_325 ? 1'h0 : _GEN_959; // @[Conditional.scala 40:58]
  assign _GEN_1020 = _T_325 ? 1'h0 : _GEN_964; // @[Conditional.scala 40:58]
  assign _GEN_1028 = io_we_i ? _GEN_972 : mstatus_spp; // @[CSR.scala 561:34]
  assign _GEN_1043 = io_we_i ? _GEN_987 : mepc_addr; // @[CSR.scala 561:34]
  assign _GEN_1044 = io_we_i ? _GEN_988 : mtvec_addr; // @[CSR.scala 561:34]
  assign _GEN_1045 = io_we_i ? _GEN_989 : medeleg; // @[CSR.scala 561:34]
  assign _GEN_1046 = io_we_i ? _GEN_990 : mideleg; // @[CSR.scala 561:34]
  assign _GEN_1048 = io_we_i ? _GEN_992 : mcause_code; // @[CSR.scala 561:34]
  assign _GEN_1050 = io_we_i ? _GEN_994 : stvec_addr; // @[CSR.scala 561:34]
  assign _GEN_1052 = io_we_i ? _GEN_996 : sepc_addr; // @[CSR.scala 561:34]
  assign _GEN_1054 = io_we_i ? _GEN_998 : scause_code; // @[CSR.scala 561:34]
  assign _GEN_1056 = io_we_i ? _GEN_1000 : sptbr_ppn; // @[CSR.scala 561:34]
  assign _GEN_1057 = io_we_i ? _GEN_1001 : mtlbindex; // @[CSR.scala 561:34]
  assign _GEN_1058 = io_we_i ? _GEN_1002 : mtlbindex_update; // @[CSR.scala 561:34]
  assign _GEN_1061 = io_we_i & _GEN_1005; // @[CSR.scala 561:34]
  assign _GEN_1066 = io_we_i & _GEN_1010; // @[CSR.scala 561:34]
  assign _GEN_1071 = io_we_i & _GEN_1015; // @[CSR.scala 561:34]
  assign _GEN_1076 = io_we_i & _GEN_1020; // @[CSR.scala 561:34]
  assign _GEN_1084 = fence_i_trap ? mstatus_spp : _GEN_1028; // @[CSR.scala 559:35]
  assign _GEN_1099 = fence_i_trap ? mepc_addr : _GEN_1043; // @[CSR.scala 559:35]
  assign _GEN_1100 = fence_i_trap ? mtvec_addr : _GEN_1044; // @[CSR.scala 559:35]
  assign _GEN_1101 = fence_i_trap ? medeleg : _GEN_1045; // @[CSR.scala 559:35]
  assign _GEN_1102 = fence_i_trap ? mideleg : _GEN_1046; // @[CSR.scala 559:35]
  assign _GEN_1104 = fence_i_trap ? mcause_code : _GEN_1048; // @[CSR.scala 559:35]
  assign _GEN_1106 = fence_i_trap ? stvec_addr : _GEN_1050; // @[CSR.scala 559:35]
  assign _GEN_1108 = fence_i_trap ? sepc_addr : _GEN_1052; // @[CSR.scala 559:35]
  assign _GEN_1110 = fence_i_trap ? scause_code : _GEN_1054; // @[CSR.scala 559:35]
  assign _GEN_1112 = fence_i_trap ? sptbr_ppn : _GEN_1056; // @[CSR.scala 559:35]
  assign _GEN_1113 = fence_i_trap ? mtlbindex : _GEN_1057; // @[CSR.scala 559:35]
  assign _GEN_1114 = fence_i_trap ? mtlbindex_update : _GEN_1058; // @[CSR.scala 559:35]
  assign _GEN_1117 = fence_i_trap ? 1'h0 : _GEN_1061; // @[CSR.scala 559:35]
  assign _GEN_1122 = fence_i_trap ? 1'h0 : _GEN_1066; // @[CSR.scala 559:35]
  assign _GEN_1127 = fence_i_trap ? 1'h0 : _GEN_1071; // @[CSR.scala 559:35]
  assign _GEN_1132 = fence_i_trap ? 1'h0 : _GEN_1076; // @[CSR.scala 559:35]
  assign _GEN_1142 = eret_from_m_trap ? mstatus_spp : _GEN_1084; // @[CSR.scala 540:39]
  assign _GEN_1155 = eret_from_m_trap ? mepc_addr : _GEN_1099; // @[CSR.scala 540:39]
  assign _GEN_1156 = eret_from_m_trap ? mtvec_addr : _GEN_1100; // @[CSR.scala 540:39]
  assign _GEN_1157 = eret_from_m_trap ? medeleg : _GEN_1101; // @[CSR.scala 540:39]
  assign _GEN_1158 = eret_from_m_trap ? mideleg : _GEN_1102; // @[CSR.scala 540:39]
  assign _GEN_1160 = eret_from_m_trap ? mcause_code : _GEN_1104; // @[CSR.scala 540:39]
  assign _GEN_1162 = eret_from_m_trap ? stvec_addr : _GEN_1106; // @[CSR.scala 540:39]
  assign _GEN_1164 = eret_from_m_trap ? sepc_addr : _GEN_1108; // @[CSR.scala 540:39]
  assign _GEN_1166 = eret_from_m_trap ? scause_code : _GEN_1110; // @[CSR.scala 540:39]
  assign _GEN_1168 = eret_from_m_trap ? sptbr_ppn : _GEN_1112; // @[CSR.scala 540:39]
  assign _GEN_1169 = eret_from_m_trap ? mtlbindex : _GEN_1113; // @[CSR.scala 540:39]
  assign _GEN_1170 = eret_from_m_trap ? mtlbindex_update : _GEN_1114; // @[CSR.scala 540:39]
  assign _GEN_1173 = eret_from_m_trap ? 1'h0 : _GEN_1117; // @[CSR.scala 540:39]
  assign _GEN_1178 = eret_from_m_trap ? 1'h0 : _GEN_1122; // @[CSR.scala 540:39]
  assign _GEN_1183 = eret_from_m_trap ? 1'h0 : _GEN_1127; // @[CSR.scala 540:39]
  assign _GEN_1188 = eret_from_m_trap ? 1'h0 : _GEN_1132; // @[CSR.scala 540:39]
  assign _GEN_1192 = eret_from_s_trap ? _GEN_130 : _GEN_1142; // @[CSR.scala 527:39]
  assign _GEN_1211 = eret_from_s_trap ? mepc_addr : _GEN_1155; // @[CSR.scala 527:39]
  assign _GEN_1212 = eret_from_s_trap ? mtvec_addr : _GEN_1156; // @[CSR.scala 527:39]
  assign _GEN_1213 = eret_from_s_trap ? medeleg : _GEN_1157; // @[CSR.scala 527:39]
  assign _GEN_1214 = eret_from_s_trap ? mideleg : _GEN_1158; // @[CSR.scala 527:39]
  assign _GEN_1216 = eret_from_s_trap ? mcause_code : _GEN_1160; // @[CSR.scala 527:39]
  assign _GEN_1218 = eret_from_s_trap ? stvec_addr : _GEN_1162; // @[CSR.scala 527:39]
  assign _GEN_1220 = eret_from_s_trap ? sepc_addr : _GEN_1164; // @[CSR.scala 527:39]
  assign _GEN_1222 = eret_from_s_trap ? scause_code : _GEN_1166; // @[CSR.scala 527:39]
  assign _GEN_1224 = eret_from_s_trap ? sptbr_ppn : _GEN_1168; // @[CSR.scala 527:39]
  assign _GEN_1225 = eret_from_s_trap ? mtlbindex : _GEN_1169; // @[CSR.scala 527:39]
  assign _GEN_1226 = eret_from_s_trap ? mtlbindex_update : _GEN_1170; // @[CSR.scala 527:39]
  assign _GEN_1229 = eret_from_s_trap ? 1'h0 : _GEN_1173; // @[CSR.scala 527:39]
  assign _GEN_1234 = eret_from_s_trap ? 1'h0 : _GEN_1178; // @[CSR.scala 527:39]
  assign _GEN_1239 = eret_from_s_trap ? 1'h0 : _GEN_1183; // @[CSR.scala 527:39]
  assign _GEN_1244 = eret_from_s_trap ? 1'h0 : _GEN_1188; // @[CSR.scala 527:39]
  assign _GEN_1247 = s_trap ? io_current_inst_addr_i[31:2] : _GEN_1220; // @[CSR.scala 474:29]
  assign _GEN_1249 = s_trap ? _GEN_120 : _GEN_1216; // @[CSR.scala 474:29]
  assign _GEN_1252 = s_trap ? _GEN_57 : {{1'd0}, _GEN_1192}; // @[CSR.scala 474:29]
  assign _GEN_1271 = s_trap ? mepc_addr : _GEN_1211; // @[CSR.scala 474:29]
  assign _GEN_1272 = s_trap ? mtvec_addr : _GEN_1212; // @[CSR.scala 474:29]
  assign _GEN_1273 = s_trap ? medeleg : _GEN_1213; // @[CSR.scala 474:29]
  assign _GEN_1274 = s_trap ? mideleg : _GEN_1214; // @[CSR.scala 474:29]
  assign _GEN_1275 = s_trap ? stvec_addr : _GEN_1218; // @[CSR.scala 474:29]
  assign _GEN_1278 = s_trap ? scause_code : _GEN_1222; // @[CSR.scala 474:29]
  assign _GEN_1280 = s_trap ? sptbr_ppn : _GEN_1224; // @[CSR.scala 474:29]
  assign _GEN_1281 = s_trap ? mtlbindex : _GEN_1225; // @[CSR.scala 474:29]
  assign _GEN_1282 = s_trap ? mtlbindex_update : _GEN_1226; // @[CSR.scala 474:29]
  assign _GEN_1285 = s_trap ? 1'h0 : _GEN_1229; // @[CSR.scala 474:29]
  assign _GEN_1290 = s_trap ? 1'h0 : _GEN_1234; // @[CSR.scala 474:29]
  assign _GEN_1295 = s_trap ? 1'h0 : _GEN_1239; // @[CSR.scala 474:29]
  assign _GEN_1300 = s_trap ? 1'h0 : _GEN_1244; // @[CSR.scala 474:29]
  assign _GEN_1303 = m_trap ? io_current_inst_addr_i[31:2] : _GEN_1271; // @[CSR.scala 416:29]
  assign _GEN_1305 = m_trap ? _GEN_86 : _GEN_1249; // @[CSR.scala 416:29]
  assign _GEN_1310 = m_trap ? sepc_addr : _GEN_1247; // @[CSR.scala 416:29]
  assign _GEN_1312 = m_trap ? {{1'd0}, mstatus_spp} : _GEN_1252; // @[CSR.scala 416:29]
  assign _GEN_1328 = m_trap ? mtvec_addr : _GEN_1272; // @[CSR.scala 416:29]
  assign _GEN_1329 = m_trap ? medeleg : _GEN_1273; // @[CSR.scala 416:29]
  assign _GEN_1330 = m_trap ? mideleg : _GEN_1274; // @[CSR.scala 416:29]
  assign _GEN_1331 = m_trap ? stvec_addr : _GEN_1275; // @[CSR.scala 416:29]
  assign _GEN_1334 = m_trap ? scause_code : _GEN_1278; // @[CSR.scala 416:29]
  assign _GEN_1336 = m_trap ? sptbr_ppn : _GEN_1280; // @[CSR.scala 416:29]
  assign _GEN_1337 = m_trap ? mtlbindex : _GEN_1281; // @[CSR.scala 416:29]
  assign _GEN_1338 = m_trap ? mtlbindex_update : _GEN_1282; // @[CSR.scala 416:29]
  assign _GEN_1341 = m_trap ? 1'h0 : _GEN_1285; // @[CSR.scala 416:29]
  assign _GEN_1346 = m_trap ? 1'h0 : _GEN_1290; // @[CSR.scala 416:29]
  assign _GEN_1351 = m_trap ? 1'h0 : _GEN_1295; // @[CSR.scala 416:29]
  assign _GEN_1356 = m_trap ? 1'h0 : _GEN_1300; // @[CSR.scala 416:29]
  assign _GEN_1359 = s_intr ? io_current_inst_addr_i[31:2] : _GEN_1310; // @[CSR.scala 384:29]
  assign _GEN_1361 = s_intr ? _GEN_53 : _GEN_1334; // @[CSR.scala 384:29]
  assign _GEN_1363 = s_intr ? _GEN_57 : _GEN_1312; // @[CSR.scala 384:29]
  assign _GEN_1365 = s_intr ? mepc_addr : _GEN_1303; // @[CSR.scala 384:29]
  assign _GEN_1367 = s_intr ? mcause_code : _GEN_1305; // @[CSR.scala 384:29]
  assign _GEN_1386 = s_intr ? mtvec_addr : _GEN_1328; // @[CSR.scala 384:29]
  assign _GEN_1387 = s_intr ? medeleg : _GEN_1329; // @[CSR.scala 384:29]
  assign _GEN_1388 = s_intr ? mideleg : _GEN_1330; // @[CSR.scala 384:29]
  assign _GEN_1389 = s_intr ? stvec_addr : _GEN_1331; // @[CSR.scala 384:29]
  assign _GEN_1392 = s_intr ? sptbr_ppn : _GEN_1336; // @[CSR.scala 384:29]
  assign _GEN_1393 = s_intr ? mtlbindex : _GEN_1337; // @[CSR.scala 384:29]
  assign _GEN_1394 = s_intr ? mtlbindex_update : _GEN_1338; // @[CSR.scala 384:29]
  assign _GEN_1397 = s_intr ? 1'h0 : _GEN_1341; // @[CSR.scala 384:29]
  assign _GEN_1402 = s_intr ? 1'h0 : _GEN_1346; // @[CSR.scala 384:29]
  assign _GEN_1407 = s_intr ? 1'h0 : _GEN_1351; // @[CSR.scala 384:29]
  assign _GEN_1412 = s_intr ? 1'h0 : _GEN_1356; // @[CSR.scala 384:29]
  assign _GEN_1415 = m_intr ? io_current_inst_addr_i[31:2] : _GEN_1365; // @[CSR.scala 350:29]
  assign _GEN_1417 = m_intr ? _GEN_37 : _GEN_1367; // @[CSR.scala 350:29]
  assign _GEN_1421 = m_intr ? sepc_addr : _GEN_1359; // @[CSR.scala 350:29]
  assign _GEN_1423 = m_intr ? scause_code : _GEN_1361; // @[CSR.scala 350:29]
  assign _GEN_1425 = m_intr ? {{1'd0}, mstatus_spp} : _GEN_1363; // @[CSR.scala 350:29]
  assign _GEN_1442 = m_intr ? mtvec_addr : _GEN_1386; // @[CSR.scala 350:29]
  assign _GEN_1443 = m_intr ? medeleg : _GEN_1387; // @[CSR.scala 350:29]
  assign _GEN_1444 = m_intr ? mideleg : _GEN_1388; // @[CSR.scala 350:29]
  assign _GEN_1445 = m_intr ? stvec_addr : _GEN_1389; // @[CSR.scala 350:29]
  assign _GEN_1448 = m_intr ? sptbr_ppn : _GEN_1392; // @[CSR.scala 350:29]
  assign _GEN_1449 = m_intr ? mtlbindex : _GEN_1393; // @[CSR.scala 350:29]
  assign _GEN_1450 = m_intr ? mtlbindex_update : _GEN_1394; // @[CSR.scala 350:29]
  assign _GEN_1453 = m_intr ? 1'h0 : _GEN_1397; // @[CSR.scala 350:29]
  assign _GEN_1458 = m_intr ? 1'h0 : _GEN_1402; // @[CSR.scala 350:29]
  assign _GEN_1463 = m_intr ? 1'h0 : _GEN_1407; // @[CSR.scala 350:29]
  assign _GEN_1468 = m_intr ? 1'h0 : _GEN_1412; // @[CSR.scala 350:29]
  assign _GEN_1471 = io_not_stall_i ? _GEN_1415 : mepc_addr; // @[CSR.scala 348:25]
  assign _GEN_1473 = io_not_stall_i ? _GEN_1417 : mcause_code; // @[CSR.scala 348:25]
  assign _GEN_1477 = io_not_stall_i ? _GEN_1421 : sepc_addr; // @[CSR.scala 348:25]
  assign _GEN_1479 = io_not_stall_i ? _GEN_1423 : scause_code; // @[CSR.scala 348:25]
  assign _GEN_1481 = io_not_stall_i ? _GEN_1425 : {{1'd0}, mstatus_spp}; // @[CSR.scala 348:25]
  assign _GEN_1498 = io_not_stall_i ? _GEN_1442 : mtvec_addr; // @[CSR.scala 348:25]
  assign _GEN_1499 = io_not_stall_i ? _GEN_1443 : medeleg; // @[CSR.scala 348:25]
  assign _GEN_1500 = io_not_stall_i ? _GEN_1444 : mideleg; // @[CSR.scala 348:25]
  assign _GEN_1501 = io_not_stall_i ? _GEN_1445 : stvec_addr; // @[CSR.scala 348:25]
  assign _GEN_1504 = io_not_stall_i ? _GEN_1448 : sptbr_ppn; // @[CSR.scala 348:25]
  assign _GEN_1505 = io_not_stall_i ? _GEN_1449 : mtlbindex; // @[CSR.scala 348:25]
  assign _GEN_1506 = io_not_stall_i ? _GEN_1450 : mtlbindex_update; // @[CSR.scala 348:25]
  assign _GEN_1509 = io_not_stall_i ? _GEN_1453 : 1'h0; // @[CSR.scala 348:25]
  assign _GEN_1514 = io_not_stall_i ? _GEN_1458 : 1'h0; // @[CSR.scala 348:25]
  assign _GEN_1519 = io_not_stall_i ? _GEN_1463 : 1'h0; // @[CSR.scala 348:25]
  assign _GEN_1524 = io_not_stall_i ? _GEN_1468 : 1'h0; // @[CSR.scala 348:25]
  assign _GEN_1527 = inst_tlb_exception ? 1'h0 : _GEN_1506; // @[CSR.scala 754:41]
  assign _GEN_1528 = inst_tlb_update ? inst_tlb_index : _GEN_1505; // @[CSR.scala 751:38]
  assign _GEN_1529 = inst_tlb_update | _GEN_1527; // @[CSR.scala 751:38]
  assign _GEN_1530 = data_tlb_exception ? 1'h0 : _GEN_1529; // @[CSR.scala 749:41]
  assign _GEN_1531 = data_tlb_exception ? _GEN_1505 : _GEN_1528; // @[CSR.scala 749:41]
  assign _GEN_1532 = data_tlb_update ? data_tlb_index : _GEN_1531; // @[CSR.scala 746:32]
  assign _GEN_1533 = data_tlb_update | _GEN_1530; // @[CSR.scala 746:32]
  assign _GEN_1539 = io_rst_n ? _GEN_1481 : 2'h0; // @[CSR.scala 283:32]
  assign _GEN_1554 = io_rst_n ? {{2'd0}, _GEN_1471} : 32'h0; // @[CSR.scala 283:32]
  assign _GEN_1555 = io_rst_n ? {{2'd0}, _GEN_1498} : 32'h0; // @[CSR.scala 283:32]
  assign _GEN_1556 = io_rst_n ? {{20'd0}, _GEN_1499} : 32'h0; // @[CSR.scala 283:32]
  assign _GEN_1557 = io_rst_n ? {{20'd0}, _GEN_1500} : 32'h0; // @[CSR.scala 283:32]
  assign _GEN_1559 = io_rst_n ? {{28'd0}, _GEN_1473} : 32'h0; // @[CSR.scala 283:32]
  assign _GEN_1561 = io_rst_n ? {{2'd0}, _GEN_1501} : 32'h0; // @[CSR.scala 283:32]
  assign _GEN_1563 = io_rst_n ? {{2'd0}, _GEN_1477} : 32'h0; // @[CSR.scala 283:32]
  assign _GEN_1565 = io_rst_n ? {{28'd0}, _GEN_1479} : 32'h0; // @[CSR.scala 283:32]
  assign _GEN_1567 = io_rst_n ? {{10'd0}, _GEN_1504} : 32'h0; // @[CSR.scala 283:32]
  assign _GEN_1568 = io_rst_n ? {{28'd0}, _GEN_1532} : 32'h0; // @[CSR.scala 283:32]
  assign _T_582 = ~io_re_i & ~io_will_write_in_mem_i; // @[CSR.scala 838:40]
  assign _T_584 = io_prv_o < io_raddr_i[9:8]; // @[CSR.scala 840:23]
  assign _T_587 = io_raddr_i[11:10] == 2'h3; // @[CSR.scala 842:73]
  assign _T_588 = io_will_write_in_mem_i & _T_587; // @[CSR.scala 842:52]
  assign _T_589 = 12'h301 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_590 = 12'hf11 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_591 = 12'hf12 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_592 = 12'hf13 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_593 = 12'hf14 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_594 = 12'h300 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_595 = 12'h305 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_596 = 12'h302 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_597 = 12'h303 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_598 = 12'h304 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_599 = 12'h344 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_600 = 12'h321 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_601 = 12'h320 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_602 = 12'h340 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_603 = 12'h341 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_604 = 12'h342 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_605 = 12'h343 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_606 = 12'h100 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_607 = 12'h105 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_608 = 12'h144 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_609 = 12'h104 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_610 = 12'h140 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_611 = 12'h141 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_612 = 12'h142 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_613 = 12'h143 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_614 = 12'h180 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_615 = 12'h7c0 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_616 = 12'h7c1 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_617 = 12'h7c2 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_618 = 12'h7c3 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_619 = 12'h7c4 == io_raddr_i; // @[Conditional.scala 37:30]
  assign _T_620 = _T_589 | _T_590; // @[Conditional.scala 37:55]
  assign _T_621 = _T_620 | _T_591; // @[Conditional.scala 37:55]
  assign _T_622 = _T_621 | _T_592; // @[Conditional.scala 37:55]
  assign _T_623 = _T_622 | _T_593; // @[Conditional.scala 37:55]
  assign _T_624 = _T_623 | _T_594; // @[Conditional.scala 37:55]
  assign _T_625 = _T_624 | _T_595; // @[Conditional.scala 37:55]
  assign _T_626 = _T_625 | _T_596; // @[Conditional.scala 37:55]
  assign _T_627 = _T_626 | _T_597; // @[Conditional.scala 37:55]
  assign _T_628 = _T_627 | _T_598; // @[Conditional.scala 37:55]
  assign _T_629 = _T_628 | _T_599; // @[Conditional.scala 37:55]
  assign _T_630 = _T_629 | _T_600; // @[Conditional.scala 37:55]
  assign _T_631 = _T_630 | _T_601; // @[Conditional.scala 37:55]
  assign _T_632 = _T_631 | _T_602; // @[Conditional.scala 37:55]
  assign _T_633 = _T_632 | _T_603; // @[Conditional.scala 37:55]
  assign _T_634 = _T_633 | _T_604; // @[Conditional.scala 37:55]
  assign _T_635 = _T_634 | _T_605; // @[Conditional.scala 37:55]
  assign _T_636 = _T_635 | _T_606; // @[Conditional.scala 37:55]
  assign _T_637 = _T_636 | _T_607; // @[Conditional.scala 37:55]
  assign _T_638 = _T_637 | _T_608; // @[Conditional.scala 37:55]
  assign _T_639 = _T_638 | _T_609; // @[Conditional.scala 37:55]
  assign _T_640 = _T_639 | _T_610; // @[Conditional.scala 37:55]
  assign _T_641 = _T_640 | _T_611; // @[Conditional.scala 37:55]
  assign _T_642 = _T_641 | _T_612; // @[Conditional.scala 37:55]
  assign _T_643 = _T_642 | _T_613; // @[Conditional.scala 37:55]
  assign _T_644 = _T_643 | _T_614; // @[Conditional.scala 37:55]
  assign _T_645 = _T_644 | _T_615; // @[Conditional.scala 37:55]
  assign _T_646 = _T_645 | _T_616; // @[Conditional.scala 37:55]
  assign _T_647 = _T_646 | _T_617; // @[Conditional.scala 37:55]
  assign _T_648 = _T_647 | _T_618; // @[Conditional.scala 37:55]
  assign _T_649 = _T_648 | _T_619; // @[Conditional.scala 37:55]
  assign _GEN_1611 = _T_588 | _T_649; // @[CSR.scala 842:90]
  assign _GEN_1612 = _T_584 | _GEN_1611; // @[CSR.scala 840:41]
  assign _GEN_1613 = _T_582 ? 1'h0 : _GEN_1612; // @[CSR.scala 838:89]
  assign _T_671 = {mstatus_fs,mstatus_mpp,1'h0,mstatus_spp,mstatus_mpie,1'h0,mstatus_spie,1'h0}; // @[Cat.scala 29:58]
  assign _T_675 = {mstatus_mie,1'h0,mstatus_sie,1'h0}; // @[Cat.scala 29:58]
  assign _T_676 = {mstatus_sd,2'h0,mstatus_vm,4'h0,mstatus_mxr,1'h0,mstatus_mprv,2'h0,_T_671,_T_675}; // @[Cat.scala 29:58]
  assign _T_678 = {mtvec_addr,2'h0}; // @[Cat.scala 29:58]
  assign _T_680 = {20'h0,medeleg}; // @[Cat.scala 29:58]
  assign _T_682 = {20'h0,mideleg}; // @[Cat.scala 29:58]
  assign _T_692 = {mip_meip,3'h0,mip_mtip,1'h0,mip_stip,1'h0,mip_msip,1'h0,mip_ssip,1'h0}; // @[Cat.scala 29:58]
  assign _T_693 = {20'h0,_T_692}; // @[Cat.scala 29:58]
  assign _T_703 = {mie_meie,3'h0,mie_mtie,1'h0,mie_stie,1'h0,mie_msie,1'h0,mie_ssie,1'h0}; // @[Cat.scala 29:58]
  assign _T_704 = {20'h0,_T_703}; // @[Cat.scala 29:58]
  assign _T_707 = {30'h0,mscounteren_tm,1'h0}; // @[Cat.scala 29:58]
  assign _T_710 = {30'h0,mucounteren_tm,1'h0}; // @[Cat.scala 29:58]
  assign _T_713 = {mepc_addr,2'h0}; // @[Cat.scala 29:58]
  assign _T_716 = {mcause_intr,27'h0,mcause_code}; // @[Cat.scala 29:58]
  assign _T_727 = {mstatus_sd,16'h0,mstatus_fs,4'h0,mstatus_spp,2'h0,mstatus_spie,3'h0,mstatus_sie,1'h0}; // @[Cat.scala 29:58]
  assign _T_729 = {stvec_addr,2'h0}; // @[Cat.scala 29:58]
  assign _T_734 = {25'h0,mip_stip,3'h0,mip_ssip,1'h0}; // @[Cat.scala 29:58]
  assign _T_739 = {25'h0,mie_stie,3'h0,mie_ssie,1'h0}; // @[Cat.scala 29:58]
  assign _T_742 = {sepc_addr,2'h0}; // @[Cat.scala 29:58]
  assign _T_745 = {scause_intr,27'h0,scause_code}; // @[Cat.scala 29:58]
  assign _T_748 = {9'h0,sptbr_ppn}; // @[Cat.scala 29:58]
  assign _T_751 = {mtlbindex_update,27'h0,mtlbindex}; // @[Cat.scala 29:58]
  assign _GEN_1618 = _T_619 ? mtlbptevaddr__T_759_data : 32'h0; // @[Conditional.scala 39:67]
  assign _GEN_1622 = _T_618 ? mtlbpte__T_757_data : _GEN_1618; // @[Conditional.scala 39:67]
  assign _GEN_1625 = _T_618 ? 1'h0 : _T_619; // @[Conditional.scala 39:67]
  assign _GEN_1629 = _T_617 ? mtlbmask__T_755_data : _GEN_1622; // @[Conditional.scala 39:67]
  assign _GEN_1632 = _T_617 ? 1'h0 : _T_618; // @[Conditional.scala 39:67]
  assign _GEN_1635 = _T_617 ? 1'h0 : _GEN_1625; // @[Conditional.scala 39:67]
  assign _GEN_1639 = _T_616 ? mtlbvpn__T_753_data : _GEN_1629; // @[Conditional.scala 39:67]
  assign _GEN_1642 = _T_616 ? 1'h0 : _T_617; // @[Conditional.scala 39:67]
  assign _GEN_1645 = _T_616 ? 1'h0 : _GEN_1632; // @[Conditional.scala 39:67]
  assign _GEN_1648 = _T_616 ? 1'h0 : _GEN_1635; // @[Conditional.scala 39:67]
  assign _GEN_1649 = _T_615 ? _T_751 : _GEN_1639; // @[Conditional.scala 39:67]
  assign _GEN_1652 = _T_615 ? 1'h0 : _T_616; // @[Conditional.scala 39:67]
  assign _GEN_1655 = _T_615 ? 1'h0 : _GEN_1642; // @[Conditional.scala 39:67]
  assign _GEN_1658 = _T_615 ? 1'h0 : _GEN_1645; // @[Conditional.scala 39:67]
  assign _GEN_1661 = _T_615 ? 1'h0 : _GEN_1648; // @[Conditional.scala 39:67]
  assign _GEN_1662 = _T_614 ? {{1'd0}, _T_748} : _GEN_1649; // @[Conditional.scala 39:67]
  assign _GEN_1665 = _T_614 ? 1'h0 : _GEN_1652; // @[Conditional.scala 39:67]
  assign _GEN_1668 = _T_614 ? 1'h0 : _GEN_1655; // @[Conditional.scala 39:67]
  assign _GEN_1671 = _T_614 ? 1'h0 : _GEN_1658; // @[Conditional.scala 39:67]
  assign _GEN_1674 = _T_614 ? 1'h0 : _GEN_1661; // @[Conditional.scala 39:67]
  assign _GEN_1675 = _T_613 ? sbadaddr : _GEN_1662; // @[Conditional.scala 39:67]
  assign _GEN_1678 = _T_613 ? 1'h0 : _GEN_1665; // @[Conditional.scala 39:67]
  assign _GEN_1681 = _T_613 ? 1'h0 : _GEN_1668; // @[Conditional.scala 39:67]
  assign _GEN_1684 = _T_613 ? 1'h0 : _GEN_1671; // @[Conditional.scala 39:67]
  assign _GEN_1687 = _T_613 ? 1'h0 : _GEN_1674; // @[Conditional.scala 39:67]
  assign _GEN_1688 = _T_612 ? _T_745 : _GEN_1675; // @[Conditional.scala 39:67]
  assign _GEN_1691 = _T_612 ? 1'h0 : _GEN_1678; // @[Conditional.scala 39:67]
  assign _GEN_1694 = _T_612 ? 1'h0 : _GEN_1681; // @[Conditional.scala 39:67]
  assign _GEN_1697 = _T_612 ? 1'h0 : _GEN_1684; // @[Conditional.scala 39:67]
  assign _GEN_1700 = _T_612 ? 1'h0 : _GEN_1687; // @[Conditional.scala 39:67]
  assign _GEN_1701 = _T_611 ? _T_742 : _GEN_1688; // @[Conditional.scala 39:67]
  assign _GEN_1704 = _T_611 ? 1'h0 : _GEN_1691; // @[Conditional.scala 39:67]
  assign _GEN_1707 = _T_611 ? 1'h0 : _GEN_1694; // @[Conditional.scala 39:67]
  assign _GEN_1710 = _T_611 ? 1'h0 : _GEN_1697; // @[Conditional.scala 39:67]
  assign _GEN_1713 = _T_611 ? 1'h0 : _GEN_1700; // @[Conditional.scala 39:67]
  assign _GEN_1714 = _T_610 ? sscratch : _GEN_1701; // @[Conditional.scala 39:67]
  assign _GEN_1717 = _T_610 ? 1'h0 : _GEN_1704; // @[Conditional.scala 39:67]
  assign _GEN_1720 = _T_610 ? 1'h0 : _GEN_1707; // @[Conditional.scala 39:67]
  assign _GEN_1723 = _T_610 ? 1'h0 : _GEN_1710; // @[Conditional.scala 39:67]
  assign _GEN_1726 = _T_610 ? 1'h0 : _GEN_1713; // @[Conditional.scala 39:67]
  assign _GEN_1727 = _T_609 ? {{1'd0}, _T_739} : _GEN_1714; // @[Conditional.scala 39:67]
  assign _GEN_1730 = _T_609 ? 1'h0 : _GEN_1717; // @[Conditional.scala 39:67]
  assign _GEN_1733 = _T_609 ? 1'h0 : _GEN_1720; // @[Conditional.scala 39:67]
  assign _GEN_1736 = _T_609 ? 1'h0 : _GEN_1723; // @[Conditional.scala 39:67]
  assign _GEN_1739 = _T_609 ? 1'h0 : _GEN_1726; // @[Conditional.scala 39:67]
  assign _GEN_1740 = _T_608 ? {{1'd0}, _T_734} : _GEN_1727; // @[Conditional.scala 39:67]
  assign _GEN_1743 = _T_608 ? 1'h0 : _GEN_1730; // @[Conditional.scala 39:67]
  assign _GEN_1746 = _T_608 ? 1'h0 : _GEN_1733; // @[Conditional.scala 39:67]
  assign _GEN_1749 = _T_608 ? 1'h0 : _GEN_1736; // @[Conditional.scala 39:67]
  assign _GEN_1752 = _T_608 ? 1'h0 : _GEN_1739; // @[Conditional.scala 39:67]
  assign _GEN_1753 = _T_607 ? _T_729 : _GEN_1740; // @[Conditional.scala 39:67]
  assign _GEN_1756 = _T_607 ? 1'h0 : _GEN_1743; // @[Conditional.scala 39:67]
  assign _GEN_1759 = _T_607 ? 1'h0 : _GEN_1746; // @[Conditional.scala 39:67]
  assign _GEN_1762 = _T_607 ? 1'h0 : _GEN_1749; // @[Conditional.scala 39:67]
  assign _GEN_1765 = _T_607 ? 1'h0 : _GEN_1752; // @[Conditional.scala 39:67]
  assign _GEN_1766 = _T_606 ? _T_727 : _GEN_1753; // @[Conditional.scala 39:67]
  assign _GEN_1769 = _T_606 ? 1'h0 : _GEN_1756; // @[Conditional.scala 39:67]
  assign _GEN_1772 = _T_606 ? 1'h0 : _GEN_1759; // @[Conditional.scala 39:67]
  assign _GEN_1775 = _T_606 ? 1'h0 : _GEN_1762; // @[Conditional.scala 39:67]
  assign _GEN_1778 = _T_606 ? 1'h0 : _GEN_1765; // @[Conditional.scala 39:67]
  assign _GEN_1779 = _T_605 ? mbadaddr : _GEN_1766; // @[Conditional.scala 39:67]
  assign _GEN_1782 = _T_605 ? 1'h0 : _GEN_1769; // @[Conditional.scala 39:67]
  assign _GEN_1785 = _T_605 ? 1'h0 : _GEN_1772; // @[Conditional.scala 39:67]
  assign _GEN_1788 = _T_605 ? 1'h0 : _GEN_1775; // @[Conditional.scala 39:67]
  assign _GEN_1791 = _T_605 ? 1'h0 : _GEN_1778; // @[Conditional.scala 39:67]
  assign _GEN_1792 = _T_604 ? _T_716 : _GEN_1779; // @[Conditional.scala 39:67]
  assign _GEN_1795 = _T_604 ? 1'h0 : _GEN_1782; // @[Conditional.scala 39:67]
  assign _GEN_1798 = _T_604 ? 1'h0 : _GEN_1785; // @[Conditional.scala 39:67]
  assign _GEN_1801 = _T_604 ? 1'h0 : _GEN_1788; // @[Conditional.scala 39:67]
  assign _GEN_1804 = _T_604 ? 1'h0 : _GEN_1791; // @[Conditional.scala 39:67]
  assign _GEN_1805 = _T_603 ? _T_713 : _GEN_1792; // @[Conditional.scala 39:67]
  assign _GEN_1808 = _T_603 ? 1'h0 : _GEN_1795; // @[Conditional.scala 39:67]
  assign _GEN_1811 = _T_603 ? 1'h0 : _GEN_1798; // @[Conditional.scala 39:67]
  assign _GEN_1814 = _T_603 ? 1'h0 : _GEN_1801; // @[Conditional.scala 39:67]
  assign _GEN_1817 = _T_603 ? 1'h0 : _GEN_1804; // @[Conditional.scala 39:67]
  assign _GEN_1818 = _T_602 ? mscratch : _GEN_1805; // @[Conditional.scala 39:67]
  assign _GEN_1821 = _T_602 ? 1'h0 : _GEN_1808; // @[Conditional.scala 39:67]
  assign _GEN_1824 = _T_602 ? 1'h0 : _GEN_1811; // @[Conditional.scala 39:67]
  assign _GEN_1827 = _T_602 ? 1'h0 : _GEN_1814; // @[Conditional.scala 39:67]
  assign _GEN_1830 = _T_602 ? 1'h0 : _GEN_1817; // @[Conditional.scala 39:67]
  assign _GEN_1831 = _T_601 ? _T_710 : _GEN_1818; // @[Conditional.scala 39:67]
  assign _GEN_1834 = _T_601 ? 1'h0 : _GEN_1821; // @[Conditional.scala 39:67]
  assign _GEN_1837 = _T_601 ? 1'h0 : _GEN_1824; // @[Conditional.scala 39:67]
  assign _GEN_1840 = _T_601 ? 1'h0 : _GEN_1827; // @[Conditional.scala 39:67]
  assign _GEN_1843 = _T_601 ? 1'h0 : _GEN_1830; // @[Conditional.scala 39:67]
  assign _GEN_1844 = _T_600 ? _T_707 : _GEN_1831; // @[Conditional.scala 39:67]
  assign _GEN_1847 = _T_600 ? 1'h0 : _GEN_1834; // @[Conditional.scala 39:67]
  assign _GEN_1850 = _T_600 ? 1'h0 : _GEN_1837; // @[Conditional.scala 39:67]
  assign _GEN_1853 = _T_600 ? 1'h0 : _GEN_1840; // @[Conditional.scala 39:67]
  assign _GEN_1856 = _T_600 ? 1'h0 : _GEN_1843; // @[Conditional.scala 39:67]
  assign _GEN_1857 = _T_598 ? _T_704 : _GEN_1844; // @[Conditional.scala 39:67]
  assign _GEN_1860 = _T_598 ? 1'h0 : _GEN_1847; // @[Conditional.scala 39:67]
  assign _GEN_1863 = _T_598 ? 1'h0 : _GEN_1850; // @[Conditional.scala 39:67]
  assign _GEN_1866 = _T_598 ? 1'h0 : _GEN_1853; // @[Conditional.scala 39:67]
  assign _GEN_1869 = _T_598 ? 1'h0 : _GEN_1856; // @[Conditional.scala 39:67]
  assign _GEN_1870 = _T_599 ? _T_693 : _GEN_1857; // @[Conditional.scala 39:67]
  assign _GEN_1873 = _T_599 ? 1'h0 : _GEN_1860; // @[Conditional.scala 39:67]
  assign _GEN_1876 = _T_599 ? 1'h0 : _GEN_1863; // @[Conditional.scala 39:67]
  assign _GEN_1879 = _T_599 ? 1'h0 : _GEN_1866; // @[Conditional.scala 39:67]
  assign _GEN_1882 = _T_599 ? 1'h0 : _GEN_1869; // @[Conditional.scala 39:67]
  assign _GEN_1883 = _T_597 ? _T_682 : _GEN_1870; // @[Conditional.scala 39:67]
  assign _GEN_1886 = _T_597 ? 1'h0 : _GEN_1873; // @[Conditional.scala 39:67]
  assign _GEN_1889 = _T_597 ? 1'h0 : _GEN_1876; // @[Conditional.scala 39:67]
  assign _GEN_1892 = _T_597 ? 1'h0 : _GEN_1879; // @[Conditional.scala 39:67]
  assign _GEN_1895 = _T_597 ? 1'h0 : _GEN_1882; // @[Conditional.scala 39:67]
  assign _GEN_1896 = _T_596 ? _T_680 : _GEN_1883; // @[Conditional.scala 39:67]
  assign _GEN_1899 = _T_596 ? 1'h0 : _GEN_1886; // @[Conditional.scala 39:67]
  assign _GEN_1902 = _T_596 ? 1'h0 : _GEN_1889; // @[Conditional.scala 39:67]
  assign _GEN_1905 = _T_596 ? 1'h0 : _GEN_1892; // @[Conditional.scala 39:67]
  assign _GEN_1908 = _T_596 ? 1'h0 : _GEN_1895; // @[Conditional.scala 39:67]
  assign _GEN_1909 = _T_595 ? _T_678 : _GEN_1896; // @[Conditional.scala 39:67]
  assign _GEN_1912 = _T_595 ? 1'h0 : _GEN_1899; // @[Conditional.scala 39:67]
  assign _GEN_1915 = _T_595 ? 1'h0 : _GEN_1902; // @[Conditional.scala 39:67]
  assign _GEN_1918 = _T_595 ? 1'h0 : _GEN_1905; // @[Conditional.scala 39:67]
  assign _GEN_1921 = _T_595 ? 1'h0 : _GEN_1908; // @[Conditional.scala 39:67]
  assign _GEN_1922 = _T_594 ? {{1'd0}, _T_676} : _GEN_1909; // @[Conditional.scala 39:67]
  assign _GEN_1925 = _T_594 ? 1'h0 : _GEN_1912; // @[Conditional.scala 39:67]
  assign _GEN_1928 = _T_594 ? 1'h0 : _GEN_1915; // @[Conditional.scala 39:67]
  assign _GEN_1931 = _T_594 ? 1'h0 : _GEN_1918; // @[Conditional.scala 39:67]
  assign _GEN_1934 = _T_594 ? 1'h0 : _GEN_1921; // @[Conditional.scala 39:67]
  assign _GEN_1935 = _T_593 ? 32'h0 : _GEN_1922; // @[Conditional.scala 39:67]
  assign _GEN_1938 = _T_593 ? 1'h0 : _GEN_1925; // @[Conditional.scala 39:67]
  assign _GEN_1941 = _T_593 ? 1'h0 : _GEN_1928; // @[Conditional.scala 39:67]
  assign _GEN_1944 = _T_593 ? 1'h0 : _GEN_1931; // @[Conditional.scala 39:67]
  assign _GEN_1947 = _T_593 ? 1'h0 : _GEN_1934; // @[Conditional.scala 39:67]
  assign _GEN_1948 = _T_592 ? 32'h0 : _GEN_1935; // @[Conditional.scala 39:67]
  assign _GEN_1951 = _T_592 ? 1'h0 : _GEN_1938; // @[Conditional.scala 39:67]
  assign _GEN_1954 = _T_592 ? 1'h0 : _GEN_1941; // @[Conditional.scala 39:67]
  assign _GEN_1957 = _T_592 ? 1'h0 : _GEN_1944; // @[Conditional.scala 39:67]
  assign _GEN_1960 = _T_592 ? 1'h0 : _GEN_1947; // @[Conditional.scala 39:67]
  assign _GEN_1961 = _T_591 ? 32'h0 : _GEN_1948; // @[Conditional.scala 39:67]
  assign _GEN_1964 = _T_591 ? 1'h0 : _GEN_1951; // @[Conditional.scala 39:67]
  assign _GEN_1967 = _T_591 ? 1'h0 : _GEN_1954; // @[Conditional.scala 39:67]
  assign _GEN_1970 = _T_591 ? 1'h0 : _GEN_1957; // @[Conditional.scala 39:67]
  assign _GEN_1973 = _T_591 ? 1'h0 : _GEN_1960; // @[Conditional.scala 39:67]
  assign _GEN_1974 = _T_590 ? 32'h0 : _GEN_1961; // @[Conditional.scala 39:67]
  assign _GEN_1977 = _T_590 ? 1'h0 : _GEN_1964; // @[Conditional.scala 39:67]
  assign _GEN_1980 = _T_590 ? 1'h0 : _GEN_1967; // @[Conditional.scala 39:67]
  assign _GEN_1983 = _T_590 ? 1'h0 : _GEN_1970; // @[Conditional.scala 39:67]
  assign _GEN_1986 = _T_590 ? 1'h0 : _GEN_1973; // @[Conditional.scala 39:67]
  assign _GEN_1987 = _T_589 ? 32'h40141101 : _GEN_1974; // @[Conditional.scala 40:58]
  assign _GEN_1990 = _T_589 ? 1'h0 : _GEN_1977; // @[Conditional.scala 40:58]
  assign _GEN_1993 = _T_589 ? 1'h0 : _GEN_1980; // @[Conditional.scala 40:58]
  assign _GEN_1996 = _T_589 ? 1'h0 : _GEN_1983; // @[Conditional.scala 40:58]
  assign _GEN_1999 = _T_589 ? 1'h0 : _GEN_1986; // @[Conditional.scala 40:58]
  assign _GEN_2000 = io_re_i ? _GEN_1987 : 32'h0; // @[CSR.scala 893:41]
  assign _GEN_2003 = io_re_i ? _GEN_1990 : 1'h0; // @[CSR.scala 893:41]
  assign _GEN_2006 = io_re_i ? _GEN_1993 : 1'h0; // @[CSR.scala 893:41]
  assign _GEN_2009 = io_re_i ? _GEN_1996 : 1'h0; // @[CSR.scala 893:41]
  assign _GEN_2012 = io_re_i ? _GEN_1999 : 1'h0; // @[CSR.scala 893:41]
  assign io_data_o = io_rst_n ? _GEN_2000 : 32'h0; // @[CSR.scala 892:15 CSR.scala 894:15 CSR.scala 896:15 CSR.scala 899:38 CSR.scala 900:38 CSR.scala 901:38 CSR.scala 902:38 CSR.scala 903:38 CSR.scala 906:19 CSR.scala 923:35 CSR.scala 924:35 CSR.scala 925:35 CSR.scala 928:19 CSR.scala 947:19 CSR.scala 965:40 CSR.scala 966:40 CSR.scala 967:40 CSR.scala 968:40 CSR.scala 971:19 CSR.scala 974:40 CSR.scala 977:19 CSR.scala 989:37 CSR.scala 992:19 CSR.scala 1000:19 CSR.scala 1007:37 CSR.scala 1008:37 CSR.scala 1011:19 CSR.scala 1016:38 CSR.scala 1017:38 CSR.scala 1020:19 CSR.scala 1025:45 CSR.scala 1026:45 CSR.scala 1027:45 CSR.scala 1028:45]
  assign io_protect_o = io_rst_n ? _GEN_1613 : 1'h0; // @[CSR.scala 837:18 CSR.scala 839:18 CSR.scala 841:18 CSR.scala 843:18 CSR.scala 845:18 CSR.scala 885:22]
  assign io_inst_phy_addr_o = mmu_conv0_io_phy_addr_o; // @[CSR.scala 791:22]
  assign io_inst_tlb_exception_o = inst_tlb_exception; // @[CSR.scala 232:27]
  assign io_data_phy_addr_o = mmu_conv1_io_phy_addr_o; // @[CSR.scala 826:22]
  assign io_data_tlb_exception_o = data_tlb_exception; // @[CSR.scala 231:27]
  assign io_flushreq = io_not_stall_i & _GEN_22; // @[CSR.scala 238:15 CSR.scala 245:19 CSR.scala 249:19 CSR.scala 253:19 CSR.scala 257:19 CSR.scala 261:19 CSR.scala 268:19 CSR.scala 276:19]
  assign io_exception_new_pc_o = io_not_stall_i ? _GEN_23 : 32'h0; // @[CSR.scala 239:25 CSR.scala 246:29 CSR.scala 250:29 CSR.scala 254:29 CSR.scala 258:29 CSR.scala 262:29 CSR.scala 269:29 CSR.scala 277:29]
  assign io_prv_o = io_rst_n ? next_prv : 2'h3; // @[CSR.scala 345:12 CSR.scala 758:13]
  assign mmu_conv0_io_rst_n = io_rst_n; // @[CSR.scala 764:22]
  assign mmu_conv0_io_tlb0_vpn_i = mtlbvpn__T_480_data; // @[CSR.scala 765:28]
  assign mmu_conv0_io_tlb0_mask_i = mtlbmask__T_482_data; // @[CSR.scala 765:110]
  assign mmu_conv0_io_tlb0_pte_i = mtlbpte__T_481_data; // @[CSR.scala 765:69]
  assign mmu_conv0_io_tlb1_vpn_i = mtlbvpn__T_483_data; // @[CSR.scala 766:28]
  assign mmu_conv0_io_tlb1_mask_i = mtlbmask__T_485_data; // @[CSR.scala 766:110]
  assign mmu_conv0_io_tlb1_pte_i = mtlbpte__T_484_data; // @[CSR.scala 766:69]
  assign mmu_conv0_io_tlb2_vpn_i = mtlbvpn__T_486_data; // @[CSR.scala 767:28]
  assign mmu_conv0_io_tlb2_mask_i = mtlbmask__T_488_data; // @[CSR.scala 767:110]
  assign mmu_conv0_io_tlb2_pte_i = mtlbpte__T_487_data; // @[CSR.scala 767:69]
  assign mmu_conv0_io_tlb3_vpn_i = mtlbvpn__T_489_data; // @[CSR.scala 768:28]
  assign mmu_conv0_io_tlb3_mask_i = mtlbmask__T_491_data; // @[CSR.scala 768:110]
  assign mmu_conv0_io_tlb3_pte_i = mtlbpte__T_490_data; // @[CSR.scala 768:69]
  assign mmu_conv0_io_tlb4_vpn_i = mtlbvpn__T_492_data; // @[CSR.scala 769:28]
  assign mmu_conv0_io_tlb4_mask_i = mtlbmask__T_494_data; // @[CSR.scala 769:110]
  assign mmu_conv0_io_tlb4_pte_i = mtlbpte__T_493_data; // @[CSR.scala 769:69]
  assign mmu_conv0_io_tlb5_vpn_i = mtlbvpn__T_495_data; // @[CSR.scala 770:28]
  assign mmu_conv0_io_tlb5_mask_i = mtlbmask__T_497_data; // @[CSR.scala 770:110]
  assign mmu_conv0_io_tlb5_pte_i = mtlbpte__T_496_data; // @[CSR.scala 770:69]
  assign mmu_conv0_io_tlb6_vpn_i = mtlbvpn__T_498_data; // @[CSR.scala 771:28]
  assign mmu_conv0_io_tlb6_mask_i = mtlbmask__T_500_data; // @[CSR.scala 771:110]
  assign mmu_conv0_io_tlb6_pte_i = mtlbpte__T_499_data; // @[CSR.scala 771:69]
  assign mmu_conv0_io_tlb7_vpn_i = mtlbvpn__T_501_data; // @[CSR.scala 772:28]
  assign mmu_conv0_io_tlb7_mask_i = mtlbmask__T_503_data; // @[CSR.scala 772:110]
  assign mmu_conv0_io_tlb7_pte_i = mtlbpte__T_502_data; // @[CSR.scala 772:69]
  assign mmu_conv0_io_tlb8_vpn_i = mtlbvpn__T_504_data; // @[CSR.scala 773:28]
  assign mmu_conv0_io_tlb8_mask_i = mtlbmask__T_506_data; // @[CSR.scala 773:110]
  assign mmu_conv0_io_tlb8_pte_i = mtlbpte__T_505_data; // @[CSR.scala 773:69]
  assign mmu_conv0_io_tlb9_vpn_i = mtlbvpn__T_507_data; // @[CSR.scala 774:28]
  assign mmu_conv0_io_tlb9_mask_i = mtlbmask__T_509_data; // @[CSR.scala 774:110]
  assign mmu_conv0_io_tlb9_pte_i = mtlbpte__T_508_data; // @[CSR.scala 774:69]
  assign mmu_conv0_io_tlb10_vpn_i = mtlbvpn__T_510_data; // @[CSR.scala 775:28]
  assign mmu_conv0_io_tlb10_mask_i = mtlbmask__T_512_data; // @[CSR.scala 775:111]
  assign mmu_conv0_io_tlb10_pte_i = mtlbpte__T_511_data; // @[CSR.scala 775:69]
  assign mmu_conv0_io_tlb11_vpn_i = mtlbvpn__T_513_data; // @[CSR.scala 776:28]
  assign mmu_conv0_io_tlb11_mask_i = mtlbmask__T_515_data; // @[CSR.scala 776:111]
  assign mmu_conv0_io_tlb11_pte_i = mtlbpte__T_514_data; // @[CSR.scala 776:69]
  assign mmu_conv0_io_tlb12_vpn_i = mtlbvpn__T_516_data; // @[CSR.scala 777:28]
  assign mmu_conv0_io_tlb12_mask_i = mtlbmask__T_518_data; // @[CSR.scala 777:111]
  assign mmu_conv0_io_tlb12_pte_i = mtlbpte__T_517_data; // @[CSR.scala 777:69]
  assign mmu_conv0_io_tlb13_vpn_i = mtlbvpn__T_519_data; // @[CSR.scala 778:28]
  assign mmu_conv0_io_tlb13_mask_i = mtlbmask__T_521_data; // @[CSR.scala 778:111]
  assign mmu_conv0_io_tlb13_pte_i = mtlbpte__T_520_data; // @[CSR.scala 778:69]
  assign mmu_conv0_io_tlb14_vpn_i = mtlbvpn__T_522_data; // @[CSR.scala 779:28]
  assign mmu_conv0_io_tlb14_mask_i = mtlbmask__T_524_data; // @[CSR.scala 779:111]
  assign mmu_conv0_io_tlb14_pte_i = mtlbpte__T_523_data; // @[CSR.scala 779:69]
  assign mmu_conv0_io_tlb15_vpn_i = mtlbvpn__T_525_data; // @[CSR.scala 780:28]
  assign mmu_conv0_io_tlb15_mask_i = mtlbmask__T_527_data; // @[CSR.scala 780:111]
  assign mmu_conv0_io_tlb15_pte_i = mtlbpte__T_526_data; // @[CSR.scala 780:69]
  assign mmu_conv0_io_vm_i = mstatus_vm; // @[CSR.scala 782:21]
  assign mmu_conv0_io_prv_i = next_prv; // @[CSR.scala 783:22]
  assign mmu_conv0_io_mxr_i = mstatus_mxr; // @[CSR.scala 784:22]
  assign mmu_conv0_io_ce_i = io_inst_ce_i; // @[CSR.scala 786:21]
  assign mmu_conv0_io_ex_i = 1'h1; // @[CSR.scala 787:21]
  assign mmu_conv0_io_we_i = 1'h0; // @[CSR.scala 788:21]
  assign mmu_conv0_io_vir_addr_i = io_inst_vir_addr_i; // @[CSR.scala 790:27]
  assign mmu_conv1_io_rst_n = io_rst_n; // @[CSR.scala 800:22]
  assign mmu_conv1_io_tlb0_vpn_i = mtlbvpn__T_528_data; // @[CSR.scala 801:28]
  assign mmu_conv1_io_tlb0_mask_i = mtlbmask__T_530_data; // @[CSR.scala 801:110]
  assign mmu_conv1_io_tlb0_pte_i = mtlbpte__T_529_data; // @[CSR.scala 801:69]
  assign mmu_conv1_io_tlb1_vpn_i = mtlbvpn__T_531_data; // @[CSR.scala 802:28]
  assign mmu_conv1_io_tlb1_mask_i = mtlbmask__T_533_data; // @[CSR.scala 802:110]
  assign mmu_conv1_io_tlb1_pte_i = mtlbpte__T_532_data; // @[CSR.scala 802:69]
  assign mmu_conv1_io_tlb2_vpn_i = mtlbvpn__T_534_data; // @[CSR.scala 803:28]
  assign mmu_conv1_io_tlb2_mask_i = mtlbmask__T_536_data; // @[CSR.scala 803:110]
  assign mmu_conv1_io_tlb2_pte_i = mtlbpte__T_535_data; // @[CSR.scala 803:69]
  assign mmu_conv1_io_tlb3_vpn_i = mtlbvpn__T_537_data; // @[CSR.scala 804:28]
  assign mmu_conv1_io_tlb3_mask_i = mtlbmask__T_539_data; // @[CSR.scala 804:110]
  assign mmu_conv1_io_tlb3_pte_i = mtlbpte__T_538_data; // @[CSR.scala 804:69]
  assign mmu_conv1_io_tlb4_vpn_i = mtlbvpn__T_540_data; // @[CSR.scala 805:28]
  assign mmu_conv1_io_tlb4_mask_i = mtlbmask__T_542_data; // @[CSR.scala 805:110]
  assign mmu_conv1_io_tlb4_pte_i = mtlbpte__T_541_data; // @[CSR.scala 805:69]
  assign mmu_conv1_io_tlb5_vpn_i = mtlbvpn__T_543_data; // @[CSR.scala 806:28]
  assign mmu_conv1_io_tlb5_mask_i = mtlbmask__T_545_data; // @[CSR.scala 806:110]
  assign mmu_conv1_io_tlb5_pte_i = mtlbpte__T_544_data; // @[CSR.scala 806:69]
  assign mmu_conv1_io_tlb6_vpn_i = mtlbvpn__T_546_data; // @[CSR.scala 807:28]
  assign mmu_conv1_io_tlb6_mask_i = mtlbmask__T_548_data; // @[CSR.scala 807:110]
  assign mmu_conv1_io_tlb6_pte_i = mtlbpte__T_547_data; // @[CSR.scala 807:69]
  assign mmu_conv1_io_tlb7_vpn_i = mtlbvpn__T_549_data; // @[CSR.scala 808:28]
  assign mmu_conv1_io_tlb7_mask_i = mtlbmask__T_551_data; // @[CSR.scala 808:110]
  assign mmu_conv1_io_tlb7_pte_i = mtlbpte__T_550_data; // @[CSR.scala 808:69]
  assign mmu_conv1_io_tlb8_vpn_i = mtlbvpn__T_552_data; // @[CSR.scala 809:28]
  assign mmu_conv1_io_tlb8_mask_i = mtlbmask__T_554_data; // @[CSR.scala 809:110]
  assign mmu_conv1_io_tlb8_pte_i = mtlbpte__T_553_data; // @[CSR.scala 809:69]
  assign mmu_conv1_io_tlb9_vpn_i = mtlbvpn__T_555_data; // @[CSR.scala 810:28]
  assign mmu_conv1_io_tlb9_mask_i = mtlbmask__T_557_data; // @[CSR.scala 810:110]
  assign mmu_conv1_io_tlb9_pte_i = mtlbpte__T_556_data; // @[CSR.scala 810:69]
  assign mmu_conv1_io_tlb10_vpn_i = mtlbvpn__T_558_data; // @[CSR.scala 811:28]
  assign mmu_conv1_io_tlb10_mask_i = mtlbmask__T_560_data; // @[CSR.scala 811:111]
  assign mmu_conv1_io_tlb10_pte_i = mtlbpte__T_559_data; // @[CSR.scala 811:69]
  assign mmu_conv1_io_tlb11_vpn_i = mtlbvpn__T_561_data; // @[CSR.scala 812:28]
  assign mmu_conv1_io_tlb11_mask_i = mtlbmask__T_563_data; // @[CSR.scala 812:111]
  assign mmu_conv1_io_tlb11_pte_i = mtlbpte__T_562_data; // @[CSR.scala 812:69]
  assign mmu_conv1_io_tlb12_vpn_i = mtlbvpn__T_564_data; // @[CSR.scala 813:28]
  assign mmu_conv1_io_tlb12_mask_i = mtlbmask__T_566_data; // @[CSR.scala 813:111]
  assign mmu_conv1_io_tlb12_pte_i = mtlbpte__T_565_data; // @[CSR.scala 813:69]
  assign mmu_conv1_io_tlb13_vpn_i = mtlbvpn__T_567_data; // @[CSR.scala 814:28]
  assign mmu_conv1_io_tlb13_mask_i = mtlbmask__T_569_data; // @[CSR.scala 814:111]
  assign mmu_conv1_io_tlb13_pte_i = mtlbpte__T_568_data; // @[CSR.scala 814:69]
  assign mmu_conv1_io_tlb14_vpn_i = mtlbvpn__T_570_data; // @[CSR.scala 815:28]
  assign mmu_conv1_io_tlb14_mask_i = mtlbmask__T_572_data; // @[CSR.scala 815:111]
  assign mmu_conv1_io_tlb14_pte_i = mtlbpte__T_571_data; // @[CSR.scala 815:69]
  assign mmu_conv1_io_tlb15_vpn_i = mtlbvpn__T_573_data; // @[CSR.scala 816:28]
  assign mmu_conv1_io_tlb15_mask_i = mtlbmask__T_575_data; // @[CSR.scala 816:111]
  assign mmu_conv1_io_tlb15_pte_i = mtlbpte__T_574_data; // @[CSR.scala 816:69]
  assign mmu_conv1_io_vm_i = mstatus_vm; // @[CSR.scala 818:21]
  assign mmu_conv1_io_prv_i = mstatus_mprv ? mstatus_mpp : next_prv; // @[CSR.scala 819:22]
  assign mmu_conv1_io_mxr_i = mstatus_mxr; // @[CSR.scala 820:22]
  assign mmu_conv1_io_ce_i = io_data_ce_i; // @[CSR.scala 822:21]
  assign mmu_conv1_io_ex_i = 1'h0; // @[CSR.scala 823:21]
  assign mmu_conv1_io_we_i = io_data_we_i; // @[CSR.scala 824:21]
  assign mmu_conv1_io_vir_addr_i = io_data_vir_addr_i; // @[CSR.scala 825:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mtlbvpn[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mtlbmask[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mtlbpte[initvar] = _RAND_2[31:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    mtlbptevaddr[initvar] = _RAND_3[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mstatus_vm = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  mstatus_mxr = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mstatus_mprv = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mstatus_fs = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mstatus_sd = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  mstatus_mpp = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mstatus_spp = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mstatus_mpie = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  mstatus_spie = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  mstatus_mie = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  mstatus_sie = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  mip_mtip = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  mip_stip = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  mie_mtie = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  mie_stie = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  mip_msip = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  mip_ssip = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  mie_msie = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  mie_ssie = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  mip_meip = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  mie_meie = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  mucounteren_tm = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  mscounteren_tm = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  mscratch = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  mepc_addr = _RAND_28[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  mtvec_addr = _RAND_29[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  medeleg = _RAND_30[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  mideleg = _RAND_31[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  mcause_intr = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  mcause_code = _RAND_33[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  mbadaddr = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  stvec_addr = _RAND_35[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  sscratch = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  sepc_addr = _RAND_37[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  scause_intr = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  scause_code = _RAND_39[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  sbadaddr = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  sptbr_ppn = _RAND_41[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  mtlbindex = _RAND_42[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  mtlbindex_update = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  inst_tlb_index = _RAND_44[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  inst_tlb_update = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  inst_tlb_exception = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  data_tlb_index = _RAND_47[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  data_tlb_update = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  data_tlb_exception = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  next_prv = _RAND_50[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge io_clk) begin
    if(mtlbvpn__T_192_en & mtlbvpn__T_192_mask) begin
      mtlbvpn[mtlbvpn__T_192_addr] <= mtlbvpn__T_192_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_196_en & mtlbvpn__T_196_mask) begin
      mtlbvpn[mtlbvpn__T_196_addr] <= mtlbvpn__T_196_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_200_en & mtlbvpn__T_200_mask) begin
      mtlbvpn[mtlbvpn__T_200_addr] <= mtlbvpn__T_200_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_204_en & mtlbvpn__T_204_mask) begin
      mtlbvpn[mtlbvpn__T_204_addr] <= mtlbvpn__T_204_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_208_en & mtlbvpn__T_208_mask) begin
      mtlbvpn[mtlbvpn__T_208_addr] <= mtlbvpn__T_208_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_212_en & mtlbvpn__T_212_mask) begin
      mtlbvpn[mtlbvpn__T_212_addr] <= mtlbvpn__T_212_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_216_en & mtlbvpn__T_216_mask) begin
      mtlbvpn[mtlbvpn__T_216_addr] <= mtlbvpn__T_216_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_220_en & mtlbvpn__T_220_mask) begin
      mtlbvpn[mtlbvpn__T_220_addr] <= mtlbvpn__T_220_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_224_en & mtlbvpn__T_224_mask) begin
      mtlbvpn[mtlbvpn__T_224_addr] <= mtlbvpn__T_224_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_228_en & mtlbvpn__T_228_mask) begin
      mtlbvpn[mtlbvpn__T_228_addr] <= mtlbvpn__T_228_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_232_en & mtlbvpn__T_232_mask) begin
      mtlbvpn[mtlbvpn__T_232_addr] <= mtlbvpn__T_232_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_236_en & mtlbvpn__T_236_mask) begin
      mtlbvpn[mtlbvpn__T_236_addr] <= mtlbvpn__T_236_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_240_en & mtlbvpn__T_240_mask) begin
      mtlbvpn[mtlbvpn__T_240_addr] <= mtlbvpn__T_240_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_244_en & mtlbvpn__T_244_mask) begin
      mtlbvpn[mtlbvpn__T_244_addr] <= mtlbvpn__T_244_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_248_en & mtlbvpn__T_248_mask) begin
      mtlbvpn[mtlbvpn__T_248_addr] <= mtlbvpn__T_248_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_252_en & mtlbvpn__T_252_mask) begin
      mtlbvpn[mtlbvpn__T_252_addr] <= mtlbvpn__T_252_data; // @[CSR.scala 121:26]
    end
    if(mtlbvpn__T_469_en & mtlbvpn__T_469_mask) begin
      mtlbvpn[mtlbvpn__T_469_addr] <= mtlbvpn__T_469_data; // @[CSR.scala 121:26]
    end
    if(mtlbmask__T_193_en & mtlbmask__T_193_mask) begin
      mtlbmask[mtlbmask__T_193_addr] <= mtlbmask__T_193_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_197_en & mtlbmask__T_197_mask) begin
      mtlbmask[mtlbmask__T_197_addr] <= mtlbmask__T_197_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_201_en & mtlbmask__T_201_mask) begin
      mtlbmask[mtlbmask__T_201_addr] <= mtlbmask__T_201_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_205_en & mtlbmask__T_205_mask) begin
      mtlbmask[mtlbmask__T_205_addr] <= mtlbmask__T_205_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_209_en & mtlbmask__T_209_mask) begin
      mtlbmask[mtlbmask__T_209_addr] <= mtlbmask__T_209_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_213_en & mtlbmask__T_213_mask) begin
      mtlbmask[mtlbmask__T_213_addr] <= mtlbmask__T_213_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_217_en & mtlbmask__T_217_mask) begin
      mtlbmask[mtlbmask__T_217_addr] <= mtlbmask__T_217_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_221_en & mtlbmask__T_221_mask) begin
      mtlbmask[mtlbmask__T_221_addr] <= mtlbmask__T_221_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_225_en & mtlbmask__T_225_mask) begin
      mtlbmask[mtlbmask__T_225_addr] <= mtlbmask__T_225_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_229_en & mtlbmask__T_229_mask) begin
      mtlbmask[mtlbmask__T_229_addr] <= mtlbmask__T_229_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_233_en & mtlbmask__T_233_mask) begin
      mtlbmask[mtlbmask__T_233_addr] <= mtlbmask__T_233_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_237_en & mtlbmask__T_237_mask) begin
      mtlbmask[mtlbmask__T_237_addr] <= mtlbmask__T_237_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_241_en & mtlbmask__T_241_mask) begin
      mtlbmask[mtlbmask__T_241_addr] <= mtlbmask__T_241_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_245_en & mtlbmask__T_245_mask) begin
      mtlbmask[mtlbmask__T_245_addr] <= mtlbmask__T_245_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_249_en & mtlbmask__T_249_mask) begin
      mtlbmask[mtlbmask__T_249_addr] <= mtlbmask__T_249_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_253_en & mtlbmask__T_253_mask) begin
      mtlbmask[mtlbmask__T_253_addr] <= mtlbmask__T_253_data; // @[CSR.scala 122:26]
    end
    if(mtlbmask__T_471_en & mtlbmask__T_471_mask) begin
      mtlbmask[mtlbmask__T_471_addr] <= mtlbmask__T_471_data; // @[CSR.scala 122:26]
    end
    if(mtlbpte__T_194_en & mtlbpte__T_194_mask) begin
      mtlbpte[mtlbpte__T_194_addr] <= mtlbpte__T_194_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_198_en & mtlbpte__T_198_mask) begin
      mtlbpte[mtlbpte__T_198_addr] <= mtlbpte__T_198_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_202_en & mtlbpte__T_202_mask) begin
      mtlbpte[mtlbpte__T_202_addr] <= mtlbpte__T_202_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_206_en & mtlbpte__T_206_mask) begin
      mtlbpte[mtlbpte__T_206_addr] <= mtlbpte__T_206_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_210_en & mtlbpte__T_210_mask) begin
      mtlbpte[mtlbpte__T_210_addr] <= mtlbpte__T_210_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_214_en & mtlbpte__T_214_mask) begin
      mtlbpte[mtlbpte__T_214_addr] <= mtlbpte__T_214_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_218_en & mtlbpte__T_218_mask) begin
      mtlbpte[mtlbpte__T_218_addr] <= mtlbpte__T_218_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_222_en & mtlbpte__T_222_mask) begin
      mtlbpte[mtlbpte__T_222_addr] <= mtlbpte__T_222_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_226_en & mtlbpte__T_226_mask) begin
      mtlbpte[mtlbpte__T_226_addr] <= mtlbpte__T_226_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_230_en & mtlbpte__T_230_mask) begin
      mtlbpte[mtlbpte__T_230_addr] <= mtlbpte__T_230_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_234_en & mtlbpte__T_234_mask) begin
      mtlbpte[mtlbpte__T_234_addr] <= mtlbpte__T_234_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_238_en & mtlbpte__T_238_mask) begin
      mtlbpte[mtlbpte__T_238_addr] <= mtlbpte__T_238_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_242_en & mtlbpte__T_242_mask) begin
      mtlbpte[mtlbpte__T_242_addr] <= mtlbpte__T_242_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_246_en & mtlbpte__T_246_mask) begin
      mtlbpte[mtlbpte__T_246_addr] <= mtlbpte__T_246_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_250_en & mtlbpte__T_250_mask) begin
      mtlbpte[mtlbpte__T_250_addr] <= mtlbpte__T_250_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_254_en & mtlbpte__T_254_mask) begin
      mtlbpte[mtlbpte__T_254_addr] <= mtlbpte__T_254_data; // @[CSR.scala 123:26]
    end
    if(mtlbpte__T_473_en & mtlbpte__T_473_mask) begin
      mtlbpte[mtlbpte__T_473_addr] <= mtlbpte__T_473_data; // @[CSR.scala 123:26]
    end
    if(mtlbptevaddr__T_195_en & mtlbptevaddr__T_195_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_195_addr] <= mtlbptevaddr__T_195_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_199_en & mtlbptevaddr__T_199_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_199_addr] <= mtlbptevaddr__T_199_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_203_en & mtlbptevaddr__T_203_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_203_addr] <= mtlbptevaddr__T_203_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_207_en & mtlbptevaddr__T_207_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_207_addr] <= mtlbptevaddr__T_207_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_211_en & mtlbptevaddr__T_211_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_211_addr] <= mtlbptevaddr__T_211_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_215_en & mtlbptevaddr__T_215_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_215_addr] <= mtlbptevaddr__T_215_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_219_en & mtlbptevaddr__T_219_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_219_addr] <= mtlbptevaddr__T_219_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_223_en & mtlbptevaddr__T_223_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_223_addr] <= mtlbptevaddr__T_223_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_227_en & mtlbptevaddr__T_227_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_227_addr] <= mtlbptevaddr__T_227_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_231_en & mtlbptevaddr__T_231_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_231_addr] <= mtlbptevaddr__T_231_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_235_en & mtlbptevaddr__T_235_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_235_addr] <= mtlbptevaddr__T_235_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_239_en & mtlbptevaddr__T_239_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_239_addr] <= mtlbptevaddr__T_239_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_243_en & mtlbptevaddr__T_243_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_243_addr] <= mtlbptevaddr__T_243_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_247_en & mtlbptevaddr__T_247_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_247_addr] <= mtlbptevaddr__T_247_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_251_en & mtlbptevaddr__T_251_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_251_addr] <= mtlbptevaddr__T_251_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_255_en & mtlbptevaddr__T_255_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_255_addr] <= mtlbptevaddr__T_255_data; // @[CSR.scala 124:26]
    end
    if(mtlbptevaddr__T_475_en & mtlbptevaddr__T_475_mask) begin
      mtlbptevaddr[mtlbptevaddr__T_475_addr] <= mtlbptevaddr__T_475_data; // @[CSR.scala 124:26]
    end
    if (~io_rst_n) begin
      mstatus_vm <= 5'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (_T_325) begin
                        if (_T_329) begin
                          mstatus_vm <= io_data_i[28:24];
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mstatus_mxr <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (_T_325) begin
                        mstatus_mxr <= io_data_i[19];
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mstatus_mprv <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (_T_325) begin
                        mstatus_mprv <= io_data_i[17];
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mstatus_fs <= 2'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (_T_325) begin
                        mstatus_fs <= io_data_i[14:13];
                      end else if (!(_T_351)) begin
                        if (!(_T_354)) begin
                          if (!(_T_360)) begin
                            if (!(_T_362)) begin
                              if (!(_T_364)) begin
                                if (!(_T_365)) begin
                                  if (!(_T_367)) begin
                                    if (!(_T_369)) begin
                                      if (!(_T_371)) begin
                                        if (!(_T_373)) begin
                                          if (!(_T_412)) begin
                                            if (_T_413) begin
                                              mstatus_fs <= io_data_i[14:13];
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mstatus_sd <= _T_1;
    end
    if (~io_rst_n) begin
      mstatus_mpp <= 2'h0;
    end else if (!(~io_not_stall_i)) begin
      if (m_intr) begin
        if (_T_264) begin
          mstatus_mpp <= 2'h0;
        end else if (_T_265) begin
          mstatus_mpp <= 2'h1;
        end else if (_T_266) begin
          mstatus_mpp <= 2'h3;
        end
      end else if (!(s_intr)) begin
        if (m_trap) begin
          if (_T_264) begin
            mstatus_mpp <= 2'h0;
          end else if (_T_265) begin
            mstatus_mpp <= 2'h1;
          end else if (_T_266) begin
            mstatus_mpp <= 2'h3;
          end
        end else if (!(s_trap)) begin
          if (!(eret_from_s_trap)) begin
            if (eret_from_m_trap) begin
              if (_T_185) begin
                mstatus_mpp <= 2'h0;
              end else if (_T_186) begin
                mstatus_mpp <= 2'h0;
              end else if (_T_187) begin
                mstatus_mpp <= 2'h0;
              end
            end else if (!(fence_i_trap)) begin
              if (io_we_i) begin
                if (_T_325) begin
                  if (_T_339) begin
                    mstatus_mpp <= io_data_i[12:11];
                  end
                end
              end
            end
          end
        end
      end
    end
    mstatus_spp <= _GEN_1539[0];
    if (~io_rst_n) begin
      mstatus_mpie <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (m_intr) begin
        if (_T_264) begin
          mstatus_mpie <= 1'h0;
        end else if (_T_265) begin
          mstatus_mpie <= mstatus_sie;
        end else if (_T_266) begin
          mstatus_mpie <= mstatus_mie;
        end
      end else if (!(s_intr)) begin
        if (m_trap) begin
          if (_T_264) begin
            mstatus_mpie <= 1'h0;
          end else if (_T_265) begin
            mstatus_mpie <= mstatus_sie;
          end else if (_T_266) begin
            mstatus_mpie <= mstatus_mie;
          end
        end else if (!(s_trap)) begin
          if (!(eret_from_s_trap)) begin
            if (eret_from_m_trap) begin
              mstatus_mpie <= _GEN_138;
            end else if (!(fence_i_trap)) begin
              if (io_we_i) begin
                if (_T_325) begin
                  mstatus_mpie <= io_data_i[7];
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mstatus_spie <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (s_intr) begin
          if (_T_264) begin
            mstatus_spie <= 1'h0;
          end else if (_T_265) begin
            mstatus_spie <= mstatus_sie;
          end
        end else if (!(m_trap)) begin
          if (s_trap) begin
            if (_T_264) begin
              mstatus_spie <= 1'h0;
            end else if (_T_265) begin
              mstatus_spie <= mstatus_sie;
            end
          end else if (eret_from_s_trap) begin
            mstatus_spie <= _GEN_129;
          end else if (!(eret_from_m_trap)) begin
            if (!(fence_i_trap)) begin
              if (io_we_i) begin
                if (_T_325) begin
                  mstatus_spie <= io_data_i[5];
                end else if (!(_T_351)) begin
                  if (!(_T_354)) begin
                    if (!(_T_360)) begin
                      if (!(_T_362)) begin
                        if (!(_T_364)) begin
                          if (!(_T_365)) begin
                            if (!(_T_367)) begin
                              if (!(_T_369)) begin
                                if (!(_T_371)) begin
                                  if (!(_T_373)) begin
                                    if (!(_T_412)) begin
                                      if (_T_413) begin
                                        mstatus_spie <= io_data_i[5];
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mstatus_mie <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (m_intr) begin
        mstatus_mie <= 1'h0;
      end else if (!(s_intr)) begin
        if (m_trap) begin
          mstatus_mie <= 1'h0;
        end else if (!(s_trap)) begin
          if (!(eret_from_s_trap)) begin
            if (eret_from_m_trap) begin
              if (!(_T_185)) begin
                if (_T_186) begin
                  mstatus_mie <= mstatus_mpie;
                end else if (_T_187) begin
                  mstatus_mie <= mstatus_mpie;
                end
              end
            end else if (!(fence_i_trap)) begin
              if (io_we_i) begin
                if (_T_325) begin
                  mstatus_mie <= io_data_i[3];
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mstatus_sie <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (s_intr) begin
          mstatus_sie <= 1'h0;
        end else if (!(m_trap)) begin
          if (s_trap) begin
            mstatus_sie <= 1'h0;
          end else if (eret_from_s_trap) begin
            if (!(_T_181)) begin
              if (_T_182) begin
                mstatus_sie <= mstatus_spie;
              end
            end
          end else if (!(eret_from_m_trap)) begin
            if (!(fence_i_trap)) begin
              if (io_we_i) begin
                if (_T_325) begin
                  mstatus_sie <= io_data_i[1];
                end else if (!(_T_351)) begin
                  if (!(_T_354)) begin
                    if (!(_T_360)) begin
                      if (!(_T_362)) begin
                        if (!(_T_364)) begin
                          if (!(_T_365)) begin
                            if (!(_T_367)) begin
                              if (!(_T_369)) begin
                                if (!(_T_371)) begin
                                  if (!(_T_373)) begin
                                    if (!(_T_412)) begin
                                      if (_T_413) begin
                                        mstatus_sie <= io_data_i[1];
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mip_mtip <= io_timer_int_i;
    end
    if (~io_rst_n) begin
      mip_stip <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (!(_T_325)) begin
                        if (_T_351) begin
                          mip_stip <= io_data_i[5];
                        end else if (!(_T_354)) begin
                          if (!(_T_360)) begin
                            if (!(_T_362)) begin
                              if (!(_T_364)) begin
                                if (!(_T_365)) begin
                                  if (!(_T_367)) begin
                                    if (!(_T_369)) begin
                                      if (!(_T_371)) begin
                                        if (!(_T_373)) begin
                                          if (!(_T_412)) begin
                                            if (!(_T_413)) begin
                                              if (!(_T_423)) begin
                                                if (_T_425) begin
                                                  mip_stip <= io_data_i[5];
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mie_mtie <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (!(_T_325)) begin
                        if (!(_T_351)) begin
                          if (_T_354) begin
                            mie_mtie <= io_data_i[7];
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mie_stie <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (!(_T_325)) begin
                        if (!(_T_351)) begin
                          if (_T_354) begin
                            mie_stie <= io_data_i[5];
                          end else if (!(_T_360)) begin
                            if (!(_T_362)) begin
                              if (!(_T_364)) begin
                                if (!(_T_365)) begin
                                  if (!(_T_367)) begin
                                    if (!(_T_369)) begin
                                      if (!(_T_371)) begin
                                        if (!(_T_373)) begin
                                          if (!(_T_412)) begin
                                            if (!(_T_413)) begin
                                              if (!(_T_423)) begin
                                                if (!(_T_425)) begin
                                                  if (_T_428) begin
                                                    mie_stie <= io_data_i[5];
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mip_msip <= io_software_int_i;
    end
    if (~io_rst_n) begin
      mip_ssip <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (!(_T_325)) begin
                        if (_T_351) begin
                          mip_ssip <= io_data_i[1];
                        end else if (!(_T_354)) begin
                          if (!(_T_360)) begin
                            if (!(_T_362)) begin
                              if (!(_T_364)) begin
                                if (!(_T_365)) begin
                                  if (!(_T_367)) begin
                                    if (!(_T_369)) begin
                                      if (!(_T_371)) begin
                                        if (!(_T_373)) begin
                                          if (!(_T_412)) begin
                                            if (!(_T_413)) begin
                                              if (!(_T_423)) begin
                                                if (_T_425) begin
                                                  mip_ssip <= io_data_i[1];
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mie_msie <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (!(_T_325)) begin
                        if (!(_T_351)) begin
                          if (_T_354) begin
                            mie_msie <= io_data_i[3];
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mie_ssie <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (!(_T_325)) begin
                        if (!(_T_351)) begin
                          if (_T_354) begin
                            mie_ssie <= io_data_i[1];
                          end else if (!(_T_360)) begin
                            if (!(_T_362)) begin
                              if (!(_T_364)) begin
                                if (!(_T_365)) begin
                                  if (!(_T_367)) begin
                                    if (!(_T_369)) begin
                                      if (!(_T_371)) begin
                                        if (!(_T_373)) begin
                                          if (!(_T_412)) begin
                                            if (!(_T_413)) begin
                                              if (!(_T_423)) begin
                                                if (!(_T_425)) begin
                                                  if (_T_428) begin
                                                    mie_ssie <= io_data_i[1];
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mip_meip <= io_external_int_i;
    end
    if (~io_rst_n) begin
      mie_meie <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (!(_T_325)) begin
                        if (!(_T_351)) begin
                          if (_T_354) begin
                            mie_meie <= io_data_i[11];
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mucounteren_tm <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (!(_T_325)) begin
                        if (!(_T_351)) begin
                          if (!(_T_354)) begin
                            if (!(_T_360)) begin
                              if (_T_362) begin
                                mucounteren_tm <= io_data_i[1];
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mscounteren_tm <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (!(_T_325)) begin
                        if (!(_T_351)) begin
                          if (!(_T_354)) begin
                            if (_T_360) begin
                              mscounteren_tm <= io_data_i[1];
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (~io_rst_n) begin
      mscratch <= 32'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (!(_T_325)) begin
                        if (!(_T_351)) begin
                          if (!(_T_354)) begin
                            if (!(_T_360)) begin
                              if (!(_T_362)) begin
                                if (_T_364) begin
                                  mscratch <= io_data_i;
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    mepc_addr <= _GEN_1554[29:0];
    mtvec_addr <= _GEN_1555[29:0];
    medeleg <= _GEN_1556[11:0];
    mideleg <= _GEN_1557[11:0];
    if (~io_rst_n) begin
      mcause_intr <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (m_intr) begin
        mcause_intr <= _GEN_36;
      end else if (!(s_intr)) begin
        if (m_trap) begin
          if (m_inst_misaligned_trap) begin
            mcause_intr <= 1'h0;
          end else if (m_inst_access_fault_trap) begin
            mcause_intr <= 1'h0;
          end else if (m_inst_illegal_trap) begin
            mcause_intr <= 1'h0;
          end else if (m_break_trap) begin
            mcause_intr <= 1'h0;
          end else if (m_load_misaligned_trap) begin
            mcause_intr <= 1'h0;
          end else if (m_load_access_fault_trap) begin
            mcause_intr <= 1'h0;
          end else if (m_store_misaligned_trap) begin
            mcause_intr <= 1'h0;
          end else if (m_store_access_fault_trap) begin
            mcause_intr <= 1'h0;
          end else if (m_ecall_from_u_trap) begin
            mcause_intr <= 1'h0;
          end else if (m_ecall_from_s_trap) begin
            mcause_intr <= 1'h0;
          end else if (m_ecall_from_m_trap) begin
            mcause_intr <= 1'h0;
          end
        end else if (s_trap) begin
          if (s_inst_misaligned_trap) begin
            mcause_intr <= 1'h0;
          end else if (s_inst_access_fault_trap) begin
            mcause_intr <= 1'h0;
          end else if (s_inst_illegal_trap) begin
            mcause_intr <= 1'h0;
          end else if (s_break_trap) begin
            mcause_intr <= 1'h0;
          end else if (s_load_misaligned_trap) begin
            mcause_intr <= 1'h0;
          end else if (s_load_access_fault_trap) begin
            mcause_intr <= 1'h0;
          end else if (s_store_misaligned_trap) begin
            mcause_intr <= 1'h0;
          end else if (s_store_access_fault_trap) begin
            mcause_intr <= 1'h0;
          end else if (s_ecall_from_u_trap) begin
            mcause_intr <= 1'h0;
          end else if (s_ecall_from_s_trap) begin
            mcause_intr <= 1'h0;
          end
        end else if (!(eret_from_s_trap)) begin
          if (!(eret_from_m_trap)) begin
            if (!(fence_i_trap)) begin
              if (io_we_i) begin
                if (!(_T_325)) begin
                  if (!(_T_351)) begin
                    if (!(_T_354)) begin
                      if (!(_T_360)) begin
                        if (!(_T_362)) begin
                          if (!(_T_364)) begin
                            if (!(_T_365)) begin
                              if (!(_T_367)) begin
                                if (!(_T_369)) begin
                                  if (!(_T_371)) begin
                                    if (_T_373) begin
                                      if (_T_409) begin
                                        mcause_intr <= io_data_i[31];
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    mcause_code <= _GEN_1559[3:0];
    if (~io_rst_n) begin
      mbadaddr <= 32'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (m_trap) begin
            if (m_inst_misaligned_trap) begin
              mbadaddr <= io_current_inst_addr_i;
            end else if (m_inst_access_fault_trap) begin
              mbadaddr <= io_current_inst_addr_i;
            end else if (!(m_inst_illegal_trap)) begin
              if (!(m_break_trap)) begin
                if (m_load_misaligned_trap) begin
                  mbadaddr <= io_current_data_addr_i;
                end else if (m_load_access_fault_trap) begin
                  mbadaddr <= io_current_data_addr_i;
                end else if (m_store_misaligned_trap) begin
                  mbadaddr <= io_current_data_addr_i;
                end else if (m_store_access_fault_trap) begin
                  mbadaddr <= io_current_data_addr_i;
                end
              end
            end
          end else if (s_trap) begin
            if (s_inst_misaligned_trap) begin
              mbadaddr <= io_current_inst_addr_i;
            end else if (s_inst_access_fault_trap) begin
              mbadaddr <= io_current_inst_addr_i;
            end else if (!(s_inst_illegal_trap)) begin
              if (!(s_break_trap)) begin
                if (s_load_misaligned_trap) begin
                  mbadaddr <= io_current_data_addr_i;
                end else if (s_load_access_fault_trap) begin
                  mbadaddr <= io_current_data_addr_i;
                end else if (s_store_misaligned_trap) begin
                  mbadaddr <= io_current_data_addr_i;
                end else if (s_store_access_fault_trap) begin
                  mbadaddr <= io_current_data_addr_i;
                end
              end
            end
          end else if (!(eret_from_s_trap)) begin
            if (!(eret_from_m_trap)) begin
              if (!(fence_i_trap)) begin
                if (io_we_i) begin
                  if (!(_T_325)) begin
                    if (!(_T_351)) begin
                      if (!(_T_354)) begin
                        if (!(_T_360)) begin
                          if (!(_T_362)) begin
                            if (!(_T_364)) begin
                              if (!(_T_365)) begin
                                if (!(_T_367)) begin
                                  if (!(_T_369)) begin
                                    if (!(_T_371)) begin
                                      if (!(_T_373)) begin
                                        if (_T_412) begin
                                          mbadaddr <= io_data_i;
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    stvec_addr <= _GEN_1561[29:0];
    if (~io_rst_n) begin
      sscratch <= 32'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (!(_T_325)) begin
                        if (!(_T_351)) begin
                          if (!(_T_354)) begin
                            if (!(_T_360)) begin
                              if (!(_T_362)) begin
                                if (!(_T_364)) begin
                                  if (!(_T_365)) begin
                                    if (!(_T_367)) begin
                                      if (!(_T_369)) begin
                                        if (!(_T_371)) begin
                                          if (!(_T_373)) begin
                                            if (!(_T_412)) begin
                                              if (!(_T_413)) begin
                                                if (!(_T_423)) begin
                                                  if (!(_T_425)) begin
                                                    if (!(_T_428)) begin
                                                      if (_T_431) begin
                                                        sscratch <= io_data_i;
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    sepc_addr <= _GEN_1563[29:0];
    if (~io_rst_n) begin
      scause_intr <= 1'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (s_intr) begin
          scause_intr <= _GEN_52;
        end else if (!(m_trap)) begin
          if (!(s_trap)) begin
            if (!(eret_from_s_trap)) begin
              if (!(eret_from_m_trap)) begin
                if (!(fence_i_trap)) begin
                  if (io_we_i) begin
                    if (!(_T_325)) begin
                      if (!(_T_351)) begin
                        if (!(_T_354)) begin
                          if (!(_T_360)) begin
                            if (!(_T_362)) begin
                              if (!(_T_364)) begin
                                if (!(_T_365)) begin
                                  if (!(_T_367)) begin
                                    if (!(_T_369)) begin
                                      if (!(_T_371)) begin
                                        if (!(_T_373)) begin
                                          if (!(_T_412)) begin
                                            if (!(_T_413)) begin
                                              if (!(_T_423)) begin
                                                if (!(_T_425)) begin
                                                  if (!(_T_428)) begin
                                                    if (!(_T_431)) begin
                                                      if (!(_T_432)) begin
                                                        if (_T_434) begin
                                                          if (_T_460) begin
                                                            scause_intr <= io_data_i[31];
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    scause_code <= _GEN_1565[3:0];
    if (~io_rst_n) begin
      sbadaddr <= 32'h0;
    end else if (!(~io_not_stall_i)) begin
      if (!(m_intr)) begin
        if (!(s_intr)) begin
          if (!(m_trap)) begin
            if (!(s_trap)) begin
              if (!(eret_from_s_trap)) begin
                if (!(eret_from_m_trap)) begin
                  if (!(fence_i_trap)) begin
                    if (io_we_i) begin
                      if (!(_T_325)) begin
                        if (!(_T_351)) begin
                          if (!(_T_354)) begin
                            if (!(_T_360)) begin
                              if (!(_T_362)) begin
                                if (!(_T_364)) begin
                                  if (!(_T_365)) begin
                                    if (!(_T_367)) begin
                                      if (!(_T_369)) begin
                                        if (!(_T_371)) begin
                                          if (!(_T_373)) begin
                                            if (!(_T_412)) begin
                                              if (!(_T_413)) begin
                                                if (!(_T_423)) begin
                                                  if (!(_T_425)) begin
                                                    if (!(_T_428)) begin
                                                      if (!(_T_431)) begin
                                                        if (!(_T_432)) begin
                                                          if (!(_T_434)) begin
                                                            if (_T_463) begin
                                                              sbadaddr <= io_data_i;
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    sptbr_ppn <= _GEN_1567[21:0];
    mtlbindex <= _GEN_1568[3:0];
    if (~io_rst_n) begin
      mtlbindex_update <= 1'h0;
    end else begin
      mtlbindex_update <= _GEN_1533;
    end
    inst_tlb_index <= mmu_conv0_io_hit_index_o;
    inst_tlb_update <= mmu_conv0_io_tlb_update_o;
    inst_tlb_exception <= mmu_conv0_io_tlb_exception_o;
    data_tlb_index <= mmu_conv1_io_hit_index_o;
    data_tlb_update <= mmu_conv1_io_tlb_update_o;
    data_tlb_exception <= mmu_conv1_io_tlb_exception_o;
    if (io_not_stall_i) begin
      if (m_intr) begin
        next_prv <= 2'h3;
      end else if (s_intr) begin
        next_prv <= 2'h1;
      end else if (m_trap) begin
        next_prv <= 2'h3;
      end else if (s_trap) begin
        next_prv <= 2'h1;
      end else if (eret_from_s_trap) begin
        if (_T_181) begin
          next_prv <= 2'h0;
        end else if (_T_182) begin
          next_prv <= 2'h1;
        end else begin
          next_prv <= io_prv_o;
        end
      end else if (eret_from_m_trap) begin
        if (_T_185) begin
          next_prv <= 2'h0;
        end else if (_T_186) begin
          next_prv <= 2'h1;
        end else if (_T_187) begin
          next_prv <= 2'h3;
        end else begin
          next_prv <= io_prv_o;
        end
      end else begin
        next_prv <= io_prv_o;
      end
    end else begin
      next_prv <= io_prv_o;
    end
  end
endmodule
